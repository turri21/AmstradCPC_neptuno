
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"24",x"24",x"3c",x"18"),
     1 => (x"00",x"00",x"fc",x"fc"),
     2 => (x"04",x"04",x"7c",x"7c"),
     3 => (x"00",x"00",x"08",x"0c"),
     4 => (x"54",x"54",x"5c",x"48"),
     5 => (x"00",x"00",x"20",x"74"),
     6 => (x"44",x"7f",x"3f",x"04"),
     7 => (x"00",x"00",x"00",x"44"),
     8 => (x"40",x"40",x"7c",x"3c"),
     9 => (x"00",x"00",x"7c",x"7c"),
    10 => (x"60",x"60",x"3c",x"1c"),
    11 => (x"3c",x"00",x"1c",x"3c"),
    12 => (x"60",x"30",x"60",x"7c"),
    13 => (x"44",x"00",x"3c",x"7c"),
    14 => (x"38",x"10",x"38",x"6c"),
    15 => (x"00",x"00",x"44",x"6c"),
    16 => (x"60",x"e0",x"bc",x"1c"),
    17 => (x"00",x"00",x"1c",x"3c"),
    18 => (x"5c",x"74",x"64",x"44"),
    19 => (x"00",x"00",x"44",x"4c"),
    20 => (x"77",x"3e",x"08",x"08"),
    21 => (x"00",x"00",x"41",x"41"),
    22 => (x"7f",x"7f",x"00",x"00"),
    23 => (x"00",x"00",x"00",x"00"),
    24 => (x"3e",x"77",x"41",x"41"),
    25 => (x"02",x"00",x"08",x"08"),
    26 => (x"02",x"03",x"01",x"01"),
    27 => (x"7f",x"00",x"01",x"02"),
    28 => (x"7f",x"7f",x"7f",x"7f"),
    29 => (x"08",x"00",x"7f",x"7f"),
    30 => (x"3e",x"1c",x"1c",x"08"),
    31 => (x"7f",x"7f",x"7f",x"3e"),
    32 => (x"1c",x"3e",x"3e",x"7f"),
    33 => (x"00",x"08",x"08",x"1c"),
    34 => (x"7c",x"7c",x"18",x"10"),
    35 => (x"00",x"00",x"10",x"18"),
    36 => (x"7c",x"7c",x"30",x"10"),
    37 => (x"10",x"00",x"10",x"30"),
    38 => (x"78",x"60",x"60",x"30"),
    39 => (x"42",x"00",x"06",x"1e"),
    40 => (x"3c",x"18",x"3c",x"66"),
    41 => (x"78",x"00",x"42",x"66"),
    42 => (x"c6",x"c2",x"6a",x"38"),
    43 => (x"60",x"00",x"38",x"6c"),
    44 => (x"00",x"60",x"00",x"00"),
    45 => (x"0e",x"00",x"60",x"00"),
    46 => (x"5d",x"5c",x"5b",x"5e"),
    47 => (x"4c",x"71",x"1e",x"0e"),
    48 => (x"bf",x"fe",x"f3",x"c2"),
    49 => (x"c0",x"4b",x"c0",x"4d"),
    50 => (x"02",x"ab",x"74",x"1e"),
    51 => (x"a6",x"c4",x"87",x"c7"),
    52 => (x"c5",x"78",x"c0",x"48"),
    53 => (x"48",x"a6",x"c4",x"87"),
    54 => (x"66",x"c4",x"78",x"c1"),
    55 => (x"ee",x"49",x"73",x"1e"),
    56 => (x"86",x"c8",x"87",x"df"),
    57 => (x"ef",x"49",x"e0",x"c0"),
    58 => (x"a5",x"c4",x"87",x"ef"),
    59 => (x"f0",x"49",x"6a",x"4a"),
    60 => (x"c6",x"f1",x"87",x"f0"),
    61 => (x"c1",x"85",x"cb",x"87"),
    62 => (x"ab",x"b7",x"c8",x"83"),
    63 => (x"87",x"c7",x"ff",x"04"),
    64 => (x"26",x"4d",x"26",x"26"),
    65 => (x"26",x"4b",x"26",x"4c"),
    66 => (x"4a",x"71",x"1e",x"4f"),
    67 => (x"5a",x"c2",x"f4",x"c2"),
    68 => (x"48",x"c2",x"f4",x"c2"),
    69 => (x"fe",x"49",x"78",x"c7"),
    70 => (x"4f",x"26",x"87",x"dd"),
    71 => (x"71",x"1e",x"73",x"1e"),
    72 => (x"aa",x"b7",x"c0",x"4a"),
    73 => (x"c2",x"87",x"d3",x"03"),
    74 => (x"05",x"bf",x"ed",x"d1"),
    75 => (x"4b",x"c1",x"87",x"c4"),
    76 => (x"4b",x"c0",x"87",x"c2"),
    77 => (x"5b",x"f1",x"d1",x"c2"),
    78 => (x"d1",x"c2",x"87",x"c4"),
    79 => (x"d1",x"c2",x"5a",x"f1"),
    80 => (x"c1",x"4a",x"bf",x"ed"),
    81 => (x"a2",x"c0",x"c1",x"9a"),
    82 => (x"87",x"e8",x"ec",x"49"),
    83 => (x"d1",x"c2",x"48",x"fc"),
    84 => (x"fe",x"78",x"bf",x"ed"),
    85 => (x"71",x"1e",x"87",x"ef"),
    86 => (x"1e",x"66",x"c4",x"4a"),
    87 => (x"fd",x"e9",x"49",x"72"),
    88 => (x"4f",x"26",x"26",x"87"),
    89 => (x"ed",x"d1",x"c2",x"1e"),
    90 => (x"d7",x"e6",x"49",x"bf"),
    91 => (x"f6",x"f3",x"c2",x"87"),
    92 => (x"78",x"bf",x"e8",x"48"),
    93 => (x"48",x"f2",x"f3",x"c2"),
    94 => (x"c2",x"78",x"bf",x"ec"),
    95 => (x"4a",x"bf",x"f6",x"f3"),
    96 => (x"99",x"ff",x"c3",x"49"),
    97 => (x"72",x"2a",x"b7",x"c8"),
    98 => (x"c2",x"b0",x"71",x"48"),
    99 => (x"26",x"58",x"fe",x"f3"),
   100 => (x"5b",x"5e",x"0e",x"4f"),
   101 => (x"71",x"0e",x"5d",x"5c"),
   102 => (x"87",x"c8",x"ff",x"4b"),
   103 => (x"48",x"f1",x"f3",x"c2"),
   104 => (x"49",x"73",x"50",x"c0"),
   105 => (x"70",x"87",x"fd",x"e5"),
   106 => (x"9c",x"c2",x"4c",x"49"),
   107 => (x"cb",x"49",x"ee",x"cb"),
   108 => (x"49",x"70",x"87",x"c3"),
   109 => (x"f1",x"f3",x"c2",x"4d"),
   110 => (x"c1",x"05",x"bf",x"97"),
   111 => (x"66",x"d0",x"87",x"e2"),
   112 => (x"fa",x"f3",x"c2",x"49"),
   113 => (x"d6",x"05",x"99",x"bf"),
   114 => (x"49",x"66",x"d4",x"87"),
   115 => (x"bf",x"f2",x"f3",x"c2"),
   116 => (x"87",x"cb",x"05",x"99"),
   117 => (x"cb",x"e5",x"49",x"73"),
   118 => (x"02",x"98",x"70",x"87"),
   119 => (x"c1",x"87",x"c1",x"c1"),
   120 => (x"87",x"c0",x"fe",x"4c"),
   121 => (x"d8",x"ca",x"49",x"75"),
   122 => (x"02",x"98",x"70",x"87"),
   123 => (x"f3",x"c2",x"87",x"c6"),
   124 => (x"50",x"c1",x"48",x"f1"),
   125 => (x"97",x"f1",x"f3",x"c2"),
   126 => (x"e3",x"c0",x"05",x"bf"),
   127 => (x"fa",x"f3",x"c2",x"87"),
   128 => (x"66",x"d0",x"49",x"bf"),
   129 => (x"d6",x"ff",x"05",x"99"),
   130 => (x"f2",x"f3",x"c2",x"87"),
   131 => (x"66",x"d4",x"49",x"bf"),
   132 => (x"ca",x"ff",x"05",x"99"),
   133 => (x"e4",x"49",x"73",x"87"),
   134 => (x"98",x"70",x"87",x"ca"),
   135 => (x"87",x"ff",x"fe",x"05"),
   136 => (x"dc",x"fb",x"48",x"74"),
   137 => (x"5b",x"5e",x"0e",x"87"),
   138 => (x"f4",x"0e",x"5d",x"5c"),
   139 => (x"4c",x"4d",x"c0",x"86"),
   140 => (x"c4",x"7e",x"bf",x"ec"),
   141 => (x"f3",x"c2",x"48",x"a6"),
   142 => (x"c1",x"78",x"bf",x"fe"),
   143 => (x"c7",x"1e",x"c0",x"1e"),
   144 => (x"87",x"cd",x"fd",x"49"),
   145 => (x"98",x"70",x"86",x"c8"),
   146 => (x"ff",x"87",x"cd",x"02"),
   147 => (x"87",x"cc",x"fb",x"49"),
   148 => (x"e3",x"49",x"da",x"c1"),
   149 => (x"4d",x"c1",x"87",x"ce"),
   150 => (x"97",x"f1",x"f3",x"c2"),
   151 => (x"87",x"c3",x"02",x"bf"),
   152 => (x"c2",x"87",x"ca",x"d5"),
   153 => (x"4b",x"bf",x"f6",x"f3"),
   154 => (x"bf",x"ed",x"d1",x"c2"),
   155 => (x"87",x"e9",x"c0",x"05"),
   156 => (x"e2",x"49",x"fd",x"c3"),
   157 => (x"fa",x"c3",x"87",x"ee"),
   158 => (x"87",x"e8",x"e2",x"49"),
   159 => (x"ff",x"c3",x"49",x"73"),
   160 => (x"c0",x"1e",x"71",x"99"),
   161 => (x"87",x"ce",x"fb",x"49"),
   162 => (x"b7",x"c8",x"49",x"73"),
   163 => (x"c1",x"1e",x"71",x"29"),
   164 => (x"87",x"c2",x"fb",x"49"),
   165 => (x"fa",x"c5",x"86",x"c8"),
   166 => (x"fa",x"f3",x"c2",x"87"),
   167 => (x"02",x"9b",x"4b",x"bf"),
   168 => (x"d1",x"c2",x"87",x"dd"),
   169 => (x"c7",x"49",x"bf",x"e9"),
   170 => (x"98",x"70",x"87",x"d7"),
   171 => (x"c0",x"87",x"c4",x"05"),
   172 => (x"c2",x"87",x"d2",x"4b"),
   173 => (x"fc",x"c6",x"49",x"e0"),
   174 => (x"ed",x"d1",x"c2",x"87"),
   175 => (x"c2",x"87",x"c6",x"58"),
   176 => (x"c0",x"48",x"e9",x"d1"),
   177 => (x"c2",x"49",x"73",x"78"),
   178 => (x"87",x"cd",x"05",x"99"),
   179 => (x"e1",x"49",x"eb",x"c3"),
   180 => (x"49",x"70",x"87",x"d2"),
   181 => (x"c2",x"02",x"99",x"c2"),
   182 => (x"73",x"4c",x"fb",x"87"),
   183 => (x"05",x"99",x"c1",x"49"),
   184 => (x"f4",x"c3",x"87",x"cd"),
   185 => (x"87",x"fc",x"e0",x"49"),
   186 => (x"99",x"c2",x"49",x"70"),
   187 => (x"fa",x"87",x"c2",x"02"),
   188 => (x"c8",x"49",x"73",x"4c"),
   189 => (x"87",x"cd",x"05",x"99"),
   190 => (x"e0",x"49",x"f5",x"c3"),
   191 => (x"49",x"70",x"87",x"e6"),
   192 => (x"d4",x"02",x"99",x"c2"),
   193 => (x"c2",x"f4",x"c2",x"87"),
   194 => (x"87",x"c9",x"02",x"bf"),
   195 => (x"c2",x"88",x"c1",x"48"),
   196 => (x"c2",x"58",x"c6",x"f4"),
   197 => (x"c1",x"4c",x"ff",x"87"),
   198 => (x"c4",x"49",x"73",x"4d"),
   199 => (x"87",x"ce",x"05",x"99"),
   200 => (x"ff",x"49",x"f2",x"c3"),
   201 => (x"70",x"87",x"fd",x"df"),
   202 => (x"02",x"99",x"c2",x"49"),
   203 => (x"f4",x"c2",x"87",x"db"),
   204 => (x"48",x"7e",x"bf",x"c2"),
   205 => (x"03",x"a8",x"b7",x"c7"),
   206 => (x"48",x"6e",x"87",x"cb"),
   207 => (x"f4",x"c2",x"80",x"c1"),
   208 => (x"c2",x"c0",x"58",x"c6"),
   209 => (x"c1",x"4c",x"fe",x"87"),
   210 => (x"49",x"fd",x"c3",x"4d"),
   211 => (x"87",x"d4",x"df",x"ff"),
   212 => (x"99",x"c2",x"49",x"70"),
   213 => (x"c2",x"87",x"d5",x"02"),
   214 => (x"02",x"bf",x"c2",x"f4"),
   215 => (x"c2",x"87",x"c9",x"c0"),
   216 => (x"c0",x"48",x"c2",x"f4"),
   217 => (x"87",x"c2",x"c0",x"78"),
   218 => (x"4d",x"c1",x"4c",x"fd"),
   219 => (x"ff",x"49",x"fa",x"c3"),
   220 => (x"70",x"87",x"f1",x"de"),
   221 => (x"02",x"99",x"c2",x"49"),
   222 => (x"f4",x"c2",x"87",x"d9"),
   223 => (x"c7",x"48",x"bf",x"c2"),
   224 => (x"c0",x"03",x"a8",x"b7"),
   225 => (x"f4",x"c2",x"87",x"c9"),
   226 => (x"78",x"c7",x"48",x"c2"),
   227 => (x"fc",x"87",x"c2",x"c0"),
   228 => (x"c0",x"4d",x"c1",x"4c"),
   229 => (x"c0",x"03",x"ac",x"b7"),
   230 => (x"66",x"c4",x"87",x"d1"),
   231 => (x"82",x"d8",x"c1",x"4a"),
   232 => (x"c6",x"c0",x"02",x"6a"),
   233 => (x"74",x"4b",x"6a",x"87"),
   234 => (x"c0",x"0f",x"73",x"49"),
   235 => (x"1e",x"f0",x"c3",x"1e"),
   236 => (x"f7",x"49",x"da",x"c1"),
   237 => (x"86",x"c8",x"87",x"db"),
   238 => (x"c0",x"02",x"98",x"70"),
   239 => (x"a6",x"c8",x"87",x"e2"),
   240 => (x"c2",x"f4",x"c2",x"48"),
   241 => (x"66",x"c8",x"78",x"bf"),
   242 => (x"c4",x"91",x"cb",x"49"),
   243 => (x"80",x"71",x"48",x"66"),
   244 => (x"bf",x"6e",x"7e",x"70"),
   245 => (x"87",x"c8",x"c0",x"02"),
   246 => (x"c8",x"4b",x"bf",x"6e"),
   247 => (x"0f",x"73",x"49",x"66"),
   248 => (x"c0",x"02",x"9d",x"75"),
   249 => (x"f4",x"c2",x"87",x"c8"),
   250 => (x"f3",x"49",x"bf",x"c2"),
   251 => (x"d1",x"c2",x"87",x"c9"),
   252 => (x"c0",x"02",x"bf",x"f1"),
   253 => (x"c2",x"49",x"87",x"dd"),
   254 => (x"98",x"70",x"87",x"c7"),
   255 => (x"87",x"d3",x"c0",x"02"),
   256 => (x"bf",x"c2",x"f4",x"c2"),
   257 => (x"87",x"ef",x"f2",x"49"),
   258 => (x"cf",x"f4",x"49",x"c0"),
   259 => (x"f1",x"d1",x"c2",x"87"),
   260 => (x"f4",x"78",x"c0",x"48"),
   261 => (x"87",x"e9",x"f3",x"8e"),
   262 => (x"5c",x"5b",x"5e",x"0e"),
   263 => (x"71",x"1e",x"0e",x"5d"),
   264 => (x"fe",x"f3",x"c2",x"4c"),
   265 => (x"cd",x"c1",x"49",x"bf"),
   266 => (x"d1",x"c1",x"4d",x"a1"),
   267 => (x"74",x"7e",x"69",x"81"),
   268 => (x"87",x"cf",x"02",x"9c"),
   269 => (x"74",x"4b",x"a5",x"c4"),
   270 => (x"fe",x"f3",x"c2",x"7b"),
   271 => (x"c8",x"f3",x"49",x"bf"),
   272 => (x"74",x"7b",x"6e",x"87"),
   273 => (x"87",x"c4",x"05",x"9c"),
   274 => (x"87",x"c2",x"4b",x"c0"),
   275 => (x"49",x"73",x"4b",x"c1"),
   276 => (x"d4",x"87",x"c9",x"f3"),
   277 => (x"87",x"c7",x"02",x"66"),
   278 => (x"70",x"87",x"da",x"49"),
   279 => (x"c0",x"87",x"c2",x"4a"),
   280 => (x"f5",x"d1",x"c2",x"4a"),
   281 => (x"d8",x"f2",x"26",x"5a"),
   282 => (x"00",x"00",x"00",x"87"),
   283 => (x"00",x"00",x"00",x"00"),
   284 => (x"00",x"00",x"00",x"00"),
   285 => (x"4a",x"71",x"1e",x"00"),
   286 => (x"49",x"bf",x"c8",x"ff"),
   287 => (x"26",x"48",x"a1",x"72"),
   288 => (x"c8",x"ff",x"1e",x"4f"),
   289 => (x"c0",x"fe",x"89",x"bf"),
   290 => (x"c0",x"c0",x"c0",x"c0"),
   291 => (x"87",x"c4",x"01",x"a9"),
   292 => (x"87",x"c2",x"4a",x"c0"),
   293 => (x"48",x"72",x"4a",x"c1"),
   294 => (x"5e",x"0e",x"4f",x"26"),
   295 => (x"0e",x"5d",x"5c",x"5b"),
   296 => (x"d4",x"ff",x"4b",x"71"),
   297 => (x"48",x"66",x"d0",x"4c"),
   298 => (x"49",x"d6",x"78",x"c0"),
   299 => (x"87",x"f4",x"db",x"ff"),
   300 => (x"6c",x"7c",x"ff",x"c3"),
   301 => (x"99",x"ff",x"c3",x"49"),
   302 => (x"c3",x"49",x"4d",x"71"),
   303 => (x"e0",x"c1",x"99",x"f0"),
   304 => (x"87",x"cb",x"05",x"a9"),
   305 => (x"6c",x"7c",x"ff",x"c3"),
   306 => (x"d0",x"98",x"c3",x"48"),
   307 => (x"c3",x"78",x"08",x"66"),
   308 => (x"4a",x"6c",x"7c",x"ff"),
   309 => (x"c3",x"31",x"c8",x"49"),
   310 => (x"4a",x"6c",x"7c",x"ff"),
   311 => (x"49",x"72",x"b2",x"71"),
   312 => (x"ff",x"c3",x"31",x"c8"),
   313 => (x"71",x"4a",x"6c",x"7c"),
   314 => (x"c8",x"49",x"72",x"b2"),
   315 => (x"7c",x"ff",x"c3",x"31"),
   316 => (x"b2",x"71",x"4a",x"6c"),
   317 => (x"c0",x"48",x"d0",x"ff"),
   318 => (x"9b",x"73",x"78",x"e0"),
   319 => (x"72",x"87",x"c2",x"02"),
   320 => (x"26",x"48",x"75",x"7b"),
   321 => (x"26",x"4c",x"26",x"4d"),
   322 => (x"1e",x"4f",x"26",x"4b"),
   323 => (x"86",x"f8",x"1e",x"73"),
   324 => (x"a6",x"c8",x"1e",x"76"),
   325 => (x"87",x"c2",x"fe",x"49"),
   326 => (x"4b",x"70",x"86",x"c4"),
   327 => (x"a8",x"c4",x"48",x"6e"),
   328 => (x"87",x"ef",x"c2",x"03"),
   329 => (x"f0",x"c3",x"4a",x"73"),
   330 => (x"aa",x"d0",x"c1",x"9a"),
   331 => (x"c1",x"87",x"c7",x"02"),
   332 => (x"c2",x"05",x"aa",x"e0"),
   333 => (x"9b",x"c3",x"87",x"dd"),
   334 => (x"c4",x"87",x"d8",x"02"),
   335 => (x"31",x"c9",x"49",x"66"),
   336 => (x"66",x"c4",x"1e",x"71"),
   337 => (x"c2",x"92",x"d4",x"4a"),
   338 => (x"72",x"49",x"c6",x"f4"),
   339 => (x"ee",x"d1",x"fe",x"81"),
   340 => (x"c2",x"86",x"c4",x"87"),
   341 => (x"f6",x"c0",x"05",x"ab"),
   342 => (x"1e",x"49",x"6e",x"87"),
   343 => (x"ff",x"49",x"e3",x"c0"),
   344 => (x"d8",x"87",x"e6",x"d9"),
   345 => (x"fb",x"d8",x"ff",x"49"),
   346 => (x"1e",x"c0",x"c8",x"87"),
   347 => (x"49",x"f6",x"e2",x"c2"),
   348 => (x"87",x"fc",x"ed",x"fd"),
   349 => (x"c0",x"48",x"d0",x"ff"),
   350 => (x"e2",x"c2",x"78",x"e0"),
   351 => (x"66",x"cc",x"1e",x"f6"),
   352 => (x"c2",x"92",x"d4",x"4a"),
   353 => (x"72",x"49",x"c6",x"f4"),
   354 => (x"ef",x"cf",x"fe",x"81"),
   355 => (x"c1",x"86",x"cc",x"87"),
   356 => (x"fe",x"c0",x"05",x"ab"),
   357 => (x"49",x"f2",x"c1",x"87"),
   358 => (x"87",x"f3",x"ea",x"fd"),
   359 => (x"1e",x"f6",x"e2",x"c2"),
   360 => (x"d4",x"4a",x"66",x"c4"),
   361 => (x"c6",x"f4",x"c2",x"92"),
   362 => (x"fe",x"81",x"72",x"49"),
   363 => (x"c4",x"87",x"ca",x"ce"),
   364 => (x"c0",x"1e",x"49",x"66"),
   365 => (x"d8",x"ff",x"49",x"e3"),
   366 => (x"49",x"d7",x"87",x"cf"),
   367 => (x"87",x"e4",x"d7",x"ff"),
   368 => (x"c2",x"1e",x"c0",x"c8"),
   369 => (x"fd",x"49",x"f6",x"e2"),
   370 => (x"cc",x"87",x"d4",x"ec"),
   371 => (x"48",x"d0",x"ff",x"86"),
   372 => (x"f8",x"78",x"e0",x"c0"),
   373 => (x"87",x"ef",x"fc",x"8e"),
   374 => (x"5c",x"5b",x"5e",x"0e"),
   375 => (x"71",x"1e",x"0e",x"5d"),
   376 => (x"4c",x"d4",x"ff",x"4d"),
   377 => (x"48",x"7e",x"66",x"d4"),
   378 => (x"06",x"a8",x"b7",x"c4"),
   379 => (x"48",x"c0",x"87",x"c5"),
   380 => (x"75",x"87",x"e6",x"c1"),
   381 => (x"d7",x"de",x"fe",x"49"),
   382 => (x"c4",x"1e",x"75",x"87"),
   383 => (x"93",x"d4",x"4b",x"66"),
   384 => (x"83",x"c6",x"f4",x"c2"),
   385 => (x"c9",x"fe",x"49",x"73"),
   386 => (x"83",x"c8",x"87",x"d3"),
   387 => (x"d0",x"ff",x"4b",x"6b"),
   388 => (x"78",x"e1",x"c8",x"48"),
   389 => (x"48",x"73",x"7c",x"dd"),
   390 => (x"70",x"98",x"ff",x"c3"),
   391 => (x"c8",x"49",x"73",x"7c"),
   392 => (x"c3",x"48",x"71",x"29"),
   393 => (x"7c",x"70",x"98",x"ff"),
   394 => (x"29",x"d0",x"49",x"73"),
   395 => (x"ff",x"c3",x"48",x"71"),
   396 => (x"73",x"7c",x"70",x"98"),
   397 => (x"70",x"28",x"d8",x"48"),
   398 => (x"7c",x"7c",x"c0",x"7c"),
   399 => (x"7c",x"7c",x"7c",x"7c"),
   400 => (x"7c",x"7c",x"7c",x"7c"),
   401 => (x"d0",x"ff",x"7c",x"7c"),
   402 => (x"78",x"e0",x"c0",x"48"),
   403 => (x"dc",x"1e",x"66",x"c4"),
   404 => (x"f4",x"d5",x"ff",x"49"),
   405 => (x"73",x"86",x"c8",x"87"),
   406 => (x"e6",x"fa",x"26",x"48"),
   407 => (x"5b",x"5e",x"0e",x"87"),
   408 => (x"1e",x"0e",x"5d",x"5c"),
   409 => (x"d4",x"ff",x"7e",x"71"),
   410 => (x"c2",x"1e",x"6e",x"4b"),
   411 => (x"fe",x"49",x"d6",x"f5"),
   412 => (x"c4",x"87",x"ea",x"c7"),
   413 => (x"9d",x"4d",x"70",x"86"),
   414 => (x"87",x"c3",x"c3",x"02"),
   415 => (x"bf",x"de",x"f5",x"c2"),
   416 => (x"fe",x"49",x"6e",x"4c"),
   417 => (x"ff",x"87",x"c9",x"dc"),
   418 => (x"c5",x"c8",x"48",x"d0"),
   419 => (x"7b",x"d6",x"c1",x"78"),
   420 => (x"7b",x"15",x"4a",x"c0"),
   421 => (x"e0",x"c0",x"82",x"c1"),
   422 => (x"f5",x"04",x"aa",x"b7"),
   423 => (x"48",x"d0",x"ff",x"87"),
   424 => (x"c5",x"c8",x"78",x"c4"),
   425 => (x"7b",x"d3",x"c1",x"78"),
   426 => (x"78",x"c4",x"7b",x"c1"),
   427 => (x"c1",x"02",x"9c",x"74"),
   428 => (x"e2",x"c2",x"87",x"fc"),
   429 => (x"c0",x"c8",x"7e",x"f6"),
   430 => (x"b7",x"c0",x"8c",x"4d"),
   431 => (x"87",x"c6",x"03",x"ac"),
   432 => (x"4d",x"a4",x"c0",x"c8"),
   433 => (x"ef",x"c2",x"4c",x"c0"),
   434 => (x"49",x"bf",x"97",x"e7"),
   435 => (x"d2",x"02",x"99",x"d0"),
   436 => (x"c2",x"1e",x"c0",x"87"),
   437 => (x"fe",x"49",x"d6",x"f5"),
   438 => (x"c4",x"87",x"de",x"c9"),
   439 => (x"4a",x"49",x"70",x"86"),
   440 => (x"c2",x"87",x"ef",x"c0"),
   441 => (x"c2",x"1e",x"f6",x"e2"),
   442 => (x"fe",x"49",x"d6",x"f5"),
   443 => (x"c4",x"87",x"ca",x"c9"),
   444 => (x"4a",x"49",x"70",x"86"),
   445 => (x"c8",x"48",x"d0",x"ff"),
   446 => (x"d4",x"c1",x"78",x"c5"),
   447 => (x"bf",x"97",x"6e",x"7b"),
   448 => (x"c1",x"48",x"6e",x"7b"),
   449 => (x"c1",x"7e",x"70",x"80"),
   450 => (x"f0",x"ff",x"05",x"8d"),
   451 => (x"48",x"d0",x"ff",x"87"),
   452 => (x"9a",x"72",x"78",x"c4"),
   453 => (x"c0",x"87",x"c5",x"05"),
   454 => (x"87",x"e5",x"c0",x"48"),
   455 => (x"f5",x"c2",x"1e",x"c1"),
   456 => (x"c6",x"fe",x"49",x"d6"),
   457 => (x"86",x"c4",x"87",x"f2"),
   458 => (x"fe",x"05",x"9c",x"74"),
   459 => (x"d0",x"ff",x"87",x"c4"),
   460 => (x"78",x"c5",x"c8",x"48"),
   461 => (x"c0",x"7b",x"d3",x"c1"),
   462 => (x"c1",x"78",x"c4",x"7b"),
   463 => (x"c0",x"87",x"c2",x"48"),
   464 => (x"4d",x"26",x"26",x"48"),
   465 => (x"4b",x"26",x"4c",x"26"),
   466 => (x"5e",x"0e",x"4f",x"26"),
   467 => (x"71",x"0e",x"5c",x"5b"),
   468 => (x"02",x"66",x"cc",x"4b"),
   469 => (x"4c",x"87",x"e8",x"c0"),
   470 => (x"02",x"8c",x"f0",x"c0"),
   471 => (x"74",x"87",x"e8",x"c0"),
   472 => (x"02",x"8a",x"c1",x"4a"),
   473 => (x"8a",x"87",x"e0",x"c0"),
   474 => (x"8a",x"87",x"dc",x"02"),
   475 => (x"c0",x"87",x"d8",x"02"),
   476 => (x"c0",x"02",x"8a",x"e0"),
   477 => (x"8a",x"c1",x"87",x"e3"),
   478 => (x"87",x"e4",x"c0",x"02"),
   479 => (x"73",x"87",x"e8",x"c0"),
   480 => (x"87",x"d9",x"fb",x"49"),
   481 => (x"74",x"87",x"e2",x"c0"),
   482 => (x"f9",x"49",x"c0",x"1e"),
   483 => (x"1e",x"74",x"87",x"ca"),
   484 => (x"c3",x"f9",x"49",x"73"),
   485 => (x"d0",x"86",x"c8",x"87"),
   486 => (x"c1",x"49",x"73",x"87"),
   487 => (x"87",x"c9",x"87",x"e9"),
   488 => (x"d5",x"c2",x"49",x"73"),
   489 => (x"c0",x"87",x"c2",x"87"),
   490 => (x"87",x"d8",x"fe",x"48"),
   491 => (x"e1",x"c2",x"1e",x"00"),
   492 => (x"c1",x"49",x"bf",x"ef"),
   493 => (x"f3",x"e1",x"c2",x"b9"),
   494 => (x"48",x"d4",x"ff",x"59"),
   495 => (x"ff",x"78",x"ff",x"c3"),
   496 => (x"e1",x"c8",x"48",x"d0"),
   497 => (x"48",x"d4",x"ff",x"78"),
   498 => (x"31",x"c4",x"78",x"c1"),
   499 => (x"d0",x"ff",x"78",x"71"),
   500 => (x"78",x"e0",x"c0",x"48"),
   501 => (x"71",x"1e",x"4f",x"26"),
   502 => (x"49",x"a2",x"c4",x"4a"),
   503 => (x"48",x"dd",x"f3",x"c2"),
   504 => (x"49",x"69",x"78",x"6a"),
   505 => (x"e1",x"c2",x"b9",x"c1"),
   506 => (x"c0",x"ff",x"59",x"f3"),
   507 => (x"c6",x"d0",x"ff",x"87"),
   508 => (x"26",x"48",x"c1",x"87"),
   509 => (x"4a",x"71",x"1e",x"4f"),
   510 => (x"c2",x"49",x"a2",x"c4"),
   511 => (x"7a",x"bf",x"dd",x"f3"),
   512 => (x"bf",x"ef",x"e1",x"c2"),
   513 => (x"1e",x"4f",x"26",x"79"),
   514 => (x"c2",x"1e",x"4a",x"71"),
   515 => (x"fe",x"49",x"d6",x"f5"),
   516 => (x"c4",x"87",x"ca",x"c1"),
   517 => (x"02",x"98",x"70",x"86"),
   518 => (x"e2",x"c2",x"87",x"dc"),
   519 => (x"f5",x"c2",x"1e",x"f6"),
   520 => (x"c4",x"fe",x"49",x"d6"),
   521 => (x"86",x"c4",x"87",x"d3"),
   522 => (x"c9",x"02",x"98",x"70"),
   523 => (x"f6",x"e2",x"c2",x"87"),
   524 => (x"87",x"e2",x"fe",x"49"),
   525 => (x"48",x"c0",x"87",x"c2"),
   526 => (x"71",x"1e",x"4f",x"26"),
   527 => (x"f5",x"c2",x"1e",x"4a"),
   528 => (x"c0",x"fe",x"49",x"d6"),
   529 => (x"86",x"c4",x"87",x"d7"),
   530 => (x"de",x"02",x"98",x"70"),
   531 => (x"f6",x"e2",x"c2",x"87"),
   532 => (x"87",x"e1",x"fe",x"49"),
   533 => (x"1e",x"f6",x"e2",x"c2"),
   534 => (x"49",x"d6",x"f5",x"c2"),
   535 => (x"87",x"dc",x"c4",x"fe"),
   536 => (x"98",x"70",x"86",x"c4"),
   537 => (x"c1",x"87",x"c4",x"02"),
   538 => (x"c0",x"87",x"c2",x"48"),
   539 => (x"00",x"4f",x"26",x"48"),
   540 => (x"1e",x"00",x"00",x"00"),
   541 => (x"bf",x"c0",x"e2",x"c2"),
   542 => (x"87",x"e1",x"f7",x"49"),
   543 => (x"4f",x"26",x"48",x"c0"),
   544 => (x"00",x"00",x"28",x"84"),
   545 => (x"54",x"53",x"4d",x"41"),
   546 => (x"20",x"44",x"41",x"52"),
   547 => (x"00",x"4d",x"4f",x"52"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

