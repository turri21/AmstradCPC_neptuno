
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"ec",x"f5",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"ec",x"f5",x"c2"),
    14 => (x"48",x"d0",x"e2",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ce",x"df"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"4a",x"71",x"86",x"fc"),
    21 => (x"69",x"49",x"c0",x"ff"),
    22 => (x"98",x"c0",x"c4",x"48"),
    23 => (x"02",x"6e",x"7e",x"70"),
    24 => (x"79",x"72",x"87",x"f5"),
    25 => (x"26",x"8e",x"fc",x"48"),
    26 => (x"1e",x"72",x"1e",x"4f"),
    27 => (x"48",x"12",x"1e",x"73"),
    28 => (x"87",x"ca",x"02",x"11"),
    29 => (x"98",x"df",x"c3",x"4b"),
    30 => (x"02",x"88",x"73",x"9b"),
    31 => (x"4b",x"26",x"87",x"f0"),
    32 => (x"4f",x"26",x"4a",x"26"),
    33 => (x"72",x"1e",x"73",x"1e"),
    34 => (x"04",x"8b",x"c1",x"1e"),
    35 => (x"48",x"12",x"87",x"ca"),
    36 => (x"87",x"c4",x"02",x"11"),
    37 => (x"87",x"f1",x"02",x"88"),
    38 => (x"4b",x"26",x"4a",x"26"),
    39 => (x"74",x"1e",x"4f",x"26"),
    40 => (x"72",x"1e",x"73",x"1e"),
    41 => (x"04",x"8b",x"c1",x"1e"),
    42 => (x"48",x"12",x"87",x"d0"),
    43 => (x"87",x"ca",x"02",x"11"),
    44 => (x"98",x"df",x"c3",x"4c"),
    45 => (x"02",x"88",x"74",x"9c"),
    46 => (x"4a",x"26",x"87",x"eb"),
    47 => (x"4c",x"26",x"4b",x"26"),
    48 => (x"73",x"1e",x"4f",x"26"),
    49 => (x"a9",x"73",x"81",x"48"),
    50 => (x"12",x"87",x"c5",x"02"),
    51 => (x"87",x"f6",x"05",x"53"),
    52 => (x"c4",x"1e",x"4f",x"26"),
    53 => (x"48",x"71",x"4a",x"66"),
    54 => (x"fb",x"05",x"51",x"12"),
    55 => (x"1e",x"4f",x"26",x"87"),
    56 => (x"11",x"4a",x"66",x"c4"),
    57 => (x"08",x"d4",x"ff",x"48"),
    58 => (x"05",x"8a",x"c1",x"78"),
    59 => (x"4f",x"26",x"87",x"f5"),
    60 => (x"4a",x"66",x"c4",x"1e"),
    61 => (x"c3",x"48",x"d4",x"ff"),
    62 => (x"51",x"68",x"78",x"ff"),
    63 => (x"f3",x"05",x"8a",x"c1"),
    64 => (x"1e",x"4f",x"26",x"87"),
    65 => (x"d4",x"ff",x"1e",x"73"),
    66 => (x"7b",x"ff",x"c3",x"4b"),
    67 => (x"ff",x"c3",x"4a",x"6b"),
    68 => (x"c8",x"49",x"6b",x"7b"),
    69 => (x"c3",x"b1",x"72",x"32"),
    70 => (x"4a",x"6b",x"7b",x"ff"),
    71 => (x"b2",x"71",x"31",x"c8"),
    72 => (x"6b",x"7b",x"ff",x"c3"),
    73 => (x"72",x"32",x"c8",x"49"),
    74 => (x"c4",x"48",x"71",x"b1"),
    75 => (x"26",x"4d",x"26",x"87"),
    76 => (x"26",x"4b",x"26",x"4c"),
    77 => (x"5b",x"5e",x"0e",x"4f"),
    78 => (x"71",x"0e",x"5d",x"5c"),
    79 => (x"4c",x"d4",x"ff",x"4a"),
    80 => (x"ff",x"c3",x"49",x"72"),
    81 => (x"c2",x"7c",x"71",x"99"),
    82 => (x"05",x"bf",x"d0",x"e2"),
    83 => (x"66",x"d0",x"87",x"c8"),
    84 => (x"d4",x"30",x"c9",x"48"),
    85 => (x"66",x"d0",x"58",x"a6"),
    86 => (x"c3",x"29",x"d8",x"49"),
    87 => (x"7c",x"71",x"99",x"ff"),
    88 => (x"d0",x"49",x"66",x"d0"),
    89 => (x"99",x"ff",x"c3",x"29"),
    90 => (x"66",x"d0",x"7c",x"71"),
    91 => (x"c3",x"29",x"c8",x"49"),
    92 => (x"7c",x"71",x"99",x"ff"),
    93 => (x"c3",x"49",x"66",x"d0"),
    94 => (x"7c",x"71",x"99",x"ff"),
    95 => (x"29",x"d0",x"49",x"72"),
    96 => (x"71",x"99",x"ff",x"c3"),
    97 => (x"c9",x"4b",x"6c",x"7c"),
    98 => (x"c3",x"4d",x"ff",x"f0"),
    99 => (x"d0",x"05",x"ab",x"ff"),
   100 => (x"7c",x"ff",x"c3",x"87"),
   101 => (x"8d",x"c1",x"4b",x"6c"),
   102 => (x"c3",x"87",x"c6",x"02"),
   103 => (x"f0",x"02",x"ab",x"ff"),
   104 => (x"fe",x"48",x"73",x"87"),
   105 => (x"c0",x"1e",x"87",x"c7"),
   106 => (x"48",x"d4",x"ff",x"49"),
   107 => (x"c1",x"78",x"ff",x"c3"),
   108 => (x"b7",x"c8",x"c3",x"81"),
   109 => (x"87",x"f1",x"04",x"a9"),
   110 => (x"73",x"1e",x"4f",x"26"),
   111 => (x"c4",x"87",x"e7",x"1e"),
   112 => (x"c0",x"4b",x"df",x"f8"),
   113 => (x"f0",x"ff",x"c0",x"1e"),
   114 => (x"fd",x"49",x"f7",x"c1"),
   115 => (x"86",x"c4",x"87",x"e7"),
   116 => (x"c0",x"05",x"a8",x"c1"),
   117 => (x"d4",x"ff",x"87",x"ea"),
   118 => (x"78",x"ff",x"c3",x"48"),
   119 => (x"c0",x"c0",x"c0",x"c1"),
   120 => (x"c0",x"1e",x"c0",x"c0"),
   121 => (x"e9",x"c1",x"f0",x"e1"),
   122 => (x"87",x"c9",x"fd",x"49"),
   123 => (x"98",x"70",x"86",x"c4"),
   124 => (x"ff",x"87",x"ca",x"05"),
   125 => (x"ff",x"c3",x"48",x"d4"),
   126 => (x"cb",x"48",x"c1",x"78"),
   127 => (x"87",x"e6",x"fe",x"87"),
   128 => (x"fe",x"05",x"8b",x"c1"),
   129 => (x"48",x"c0",x"87",x"fd"),
   130 => (x"1e",x"87",x"e6",x"fc"),
   131 => (x"d4",x"ff",x"1e",x"73"),
   132 => (x"78",x"ff",x"c3",x"48"),
   133 => (x"1e",x"c0",x"4b",x"d3"),
   134 => (x"c1",x"f0",x"ff",x"c0"),
   135 => (x"d4",x"fc",x"49",x"c1"),
   136 => (x"70",x"86",x"c4",x"87"),
   137 => (x"87",x"ca",x"05",x"98"),
   138 => (x"c3",x"48",x"d4",x"ff"),
   139 => (x"48",x"c1",x"78",x"ff"),
   140 => (x"f1",x"fd",x"87",x"cb"),
   141 => (x"05",x"8b",x"c1",x"87"),
   142 => (x"c0",x"87",x"db",x"ff"),
   143 => (x"87",x"f1",x"fb",x"48"),
   144 => (x"5c",x"5b",x"5e",x"0e"),
   145 => (x"4c",x"d4",x"ff",x"0e"),
   146 => (x"c6",x"87",x"db",x"fd"),
   147 => (x"e1",x"c0",x"1e",x"ea"),
   148 => (x"49",x"c8",x"c1",x"f0"),
   149 => (x"c4",x"87",x"de",x"fb"),
   150 => (x"02",x"a8",x"c1",x"86"),
   151 => (x"ea",x"fe",x"87",x"c8"),
   152 => (x"c1",x"48",x"c0",x"87"),
   153 => (x"da",x"fa",x"87",x"e2"),
   154 => (x"cf",x"49",x"70",x"87"),
   155 => (x"c6",x"99",x"ff",x"ff"),
   156 => (x"c8",x"02",x"a9",x"ea"),
   157 => (x"87",x"d3",x"fe",x"87"),
   158 => (x"cb",x"c1",x"48",x"c0"),
   159 => (x"7c",x"ff",x"c3",x"87"),
   160 => (x"fc",x"4b",x"f1",x"c0"),
   161 => (x"98",x"70",x"87",x"f4"),
   162 => (x"87",x"eb",x"c0",x"02"),
   163 => (x"ff",x"c0",x"1e",x"c0"),
   164 => (x"49",x"fa",x"c1",x"f0"),
   165 => (x"c4",x"87",x"de",x"fa"),
   166 => (x"05",x"98",x"70",x"86"),
   167 => (x"ff",x"c3",x"87",x"d9"),
   168 => (x"c3",x"49",x"6c",x"7c"),
   169 => (x"7c",x"7c",x"7c",x"ff"),
   170 => (x"99",x"c0",x"c1",x"7c"),
   171 => (x"c1",x"87",x"c4",x"02"),
   172 => (x"c0",x"87",x"d5",x"48"),
   173 => (x"c2",x"87",x"d1",x"48"),
   174 => (x"87",x"c4",x"05",x"ab"),
   175 => (x"87",x"c8",x"48",x"c0"),
   176 => (x"fe",x"05",x"8b",x"c1"),
   177 => (x"48",x"c0",x"87",x"fd"),
   178 => (x"1e",x"87",x"e4",x"f9"),
   179 => (x"e2",x"c2",x"1e",x"73"),
   180 => (x"78",x"c1",x"48",x"d0"),
   181 => (x"d0",x"ff",x"4b",x"c7"),
   182 => (x"fb",x"78",x"c2",x"48"),
   183 => (x"d0",x"ff",x"87",x"c8"),
   184 => (x"c0",x"78",x"c3",x"48"),
   185 => (x"d0",x"e5",x"c0",x"1e"),
   186 => (x"f9",x"49",x"c0",x"c1"),
   187 => (x"86",x"c4",x"87",x"c7"),
   188 => (x"c1",x"05",x"a8",x"c1"),
   189 => (x"ab",x"c2",x"4b",x"87"),
   190 => (x"c0",x"87",x"c5",x"05"),
   191 => (x"87",x"f9",x"c0",x"48"),
   192 => (x"ff",x"05",x"8b",x"c1"),
   193 => (x"f7",x"fc",x"87",x"d0"),
   194 => (x"d4",x"e2",x"c2",x"87"),
   195 => (x"05",x"98",x"70",x"58"),
   196 => (x"1e",x"c1",x"87",x"cd"),
   197 => (x"c1",x"f0",x"ff",x"c0"),
   198 => (x"d8",x"f8",x"49",x"d0"),
   199 => (x"ff",x"86",x"c4",x"87"),
   200 => (x"ff",x"c3",x"48",x"d4"),
   201 => (x"87",x"e0",x"c4",x"78"),
   202 => (x"58",x"d8",x"e2",x"c2"),
   203 => (x"c2",x"48",x"d0",x"ff"),
   204 => (x"48",x"d4",x"ff",x"78"),
   205 => (x"c1",x"78",x"ff",x"c3"),
   206 => (x"87",x"f5",x"f7",x"48"),
   207 => (x"5c",x"5b",x"5e",x"0e"),
   208 => (x"4a",x"71",x"0e",x"5d"),
   209 => (x"ff",x"4d",x"ff",x"c3"),
   210 => (x"7c",x"75",x"4c",x"d4"),
   211 => (x"c4",x"48",x"d0",x"ff"),
   212 => (x"7c",x"75",x"78",x"c3"),
   213 => (x"ff",x"c0",x"1e",x"72"),
   214 => (x"49",x"d8",x"c1",x"f0"),
   215 => (x"c4",x"87",x"d6",x"f7"),
   216 => (x"02",x"98",x"70",x"86"),
   217 => (x"48",x"c0",x"87",x"c5"),
   218 => (x"75",x"87",x"f0",x"c0"),
   219 => (x"7c",x"fe",x"c3",x"7c"),
   220 => (x"d4",x"1e",x"c0",x"c8"),
   221 => (x"e6",x"f5",x"49",x"66"),
   222 => (x"75",x"86",x"c4",x"87"),
   223 => (x"75",x"7c",x"75",x"7c"),
   224 => (x"e0",x"da",x"d8",x"7c"),
   225 => (x"6c",x"7c",x"75",x"4b"),
   226 => (x"c5",x"05",x"99",x"49"),
   227 => (x"05",x"8b",x"c1",x"87"),
   228 => (x"7c",x"75",x"87",x"f3"),
   229 => (x"c2",x"48",x"d0",x"ff"),
   230 => (x"f6",x"48",x"c1",x"78"),
   231 => (x"ff",x"1e",x"87",x"cf"),
   232 => (x"d0",x"ff",x"4a",x"d4"),
   233 => (x"78",x"d1",x"c4",x"48"),
   234 => (x"c1",x"7a",x"ff",x"c3"),
   235 => (x"87",x"f8",x"05",x"89"),
   236 => (x"73",x"1e",x"4f",x"26"),
   237 => (x"c5",x"4b",x"71",x"1e"),
   238 => (x"4a",x"df",x"cd",x"ee"),
   239 => (x"c3",x"48",x"d4",x"ff"),
   240 => (x"48",x"68",x"78",x"ff"),
   241 => (x"02",x"a8",x"fe",x"c3"),
   242 => (x"8a",x"c1",x"87",x"c5"),
   243 => (x"72",x"87",x"ed",x"05"),
   244 => (x"87",x"c5",x"05",x"9a"),
   245 => (x"ea",x"c0",x"48",x"c0"),
   246 => (x"02",x"9b",x"73",x"87"),
   247 => (x"66",x"c8",x"87",x"cc"),
   248 => (x"f4",x"49",x"73",x"1e"),
   249 => (x"86",x"c4",x"87",x"ca"),
   250 => (x"66",x"c8",x"87",x"c6"),
   251 => (x"87",x"ee",x"fe",x"49"),
   252 => (x"c3",x"48",x"d4",x"ff"),
   253 => (x"73",x"78",x"78",x"ff"),
   254 => (x"87",x"c5",x"05",x"9b"),
   255 => (x"d0",x"48",x"d0",x"ff"),
   256 => (x"f4",x"48",x"c1",x"78"),
   257 => (x"73",x"1e",x"87",x"eb"),
   258 => (x"c0",x"4a",x"71",x"1e"),
   259 => (x"48",x"d4",x"ff",x"4b"),
   260 => (x"ff",x"78",x"ff",x"c3"),
   261 => (x"c3",x"c4",x"48",x"d0"),
   262 => (x"48",x"d4",x"ff",x"78"),
   263 => (x"72",x"78",x"ff",x"c3"),
   264 => (x"f0",x"ff",x"c0",x"1e"),
   265 => (x"f4",x"49",x"d1",x"c1"),
   266 => (x"86",x"c4",x"87",x"cb"),
   267 => (x"cd",x"05",x"98",x"70"),
   268 => (x"1e",x"c0",x"c8",x"87"),
   269 => (x"fd",x"49",x"66",x"cc"),
   270 => (x"86",x"c4",x"87",x"f8"),
   271 => (x"d0",x"ff",x"4b",x"70"),
   272 => (x"73",x"78",x"c2",x"48"),
   273 => (x"87",x"e9",x"f3",x"48"),
   274 => (x"5c",x"5b",x"5e",x"0e"),
   275 => (x"1e",x"c0",x"0e",x"5d"),
   276 => (x"c1",x"f0",x"ff",x"c0"),
   277 => (x"dc",x"f3",x"49",x"c9"),
   278 => (x"c2",x"1e",x"d2",x"87"),
   279 => (x"fd",x"49",x"d8",x"e2"),
   280 => (x"86",x"c8",x"87",x"d0"),
   281 => (x"84",x"c1",x"4c",x"c0"),
   282 => (x"04",x"ac",x"b7",x"d2"),
   283 => (x"e2",x"c2",x"87",x"f8"),
   284 => (x"49",x"bf",x"97",x"d8"),
   285 => (x"c1",x"99",x"c0",x"c3"),
   286 => (x"c0",x"05",x"a9",x"c0"),
   287 => (x"e2",x"c2",x"87",x"e7"),
   288 => (x"49",x"bf",x"97",x"df"),
   289 => (x"e2",x"c2",x"31",x"d0"),
   290 => (x"4a",x"bf",x"97",x"e0"),
   291 => (x"b1",x"72",x"32",x"c8"),
   292 => (x"97",x"e1",x"e2",x"c2"),
   293 => (x"71",x"b1",x"4a",x"bf"),
   294 => (x"ff",x"ff",x"cf",x"4c"),
   295 => (x"84",x"c1",x"9c",x"ff"),
   296 => (x"e7",x"c1",x"34",x"ca"),
   297 => (x"e1",x"e2",x"c2",x"87"),
   298 => (x"c1",x"49",x"bf",x"97"),
   299 => (x"c2",x"99",x"c6",x"31"),
   300 => (x"bf",x"97",x"e2",x"e2"),
   301 => (x"2a",x"b7",x"c7",x"4a"),
   302 => (x"e2",x"c2",x"b1",x"72"),
   303 => (x"4a",x"bf",x"97",x"dd"),
   304 => (x"c2",x"9d",x"cf",x"4d"),
   305 => (x"bf",x"97",x"de",x"e2"),
   306 => (x"ca",x"9a",x"c3",x"4a"),
   307 => (x"df",x"e2",x"c2",x"32"),
   308 => (x"c2",x"4b",x"bf",x"97"),
   309 => (x"c2",x"b2",x"73",x"33"),
   310 => (x"bf",x"97",x"e0",x"e2"),
   311 => (x"9b",x"c0",x"c3",x"4b"),
   312 => (x"73",x"2b",x"b7",x"c6"),
   313 => (x"c1",x"81",x"c2",x"b2"),
   314 => (x"70",x"30",x"71",x"48"),
   315 => (x"75",x"48",x"c1",x"49"),
   316 => (x"72",x"4d",x"70",x"30"),
   317 => (x"71",x"84",x"c1",x"4c"),
   318 => (x"b7",x"c0",x"c8",x"94"),
   319 => (x"87",x"cc",x"06",x"ad"),
   320 => (x"2d",x"b7",x"34",x"c1"),
   321 => (x"ad",x"b7",x"c0",x"c8"),
   322 => (x"87",x"f4",x"ff",x"01"),
   323 => (x"dc",x"f0",x"48",x"74"),
   324 => (x"5b",x"5e",x"0e",x"87"),
   325 => (x"f8",x"0e",x"5d",x"5c"),
   326 => (x"fe",x"ea",x"c2",x"86"),
   327 => (x"c2",x"78",x"c0",x"48"),
   328 => (x"c0",x"1e",x"f6",x"e2"),
   329 => (x"87",x"de",x"fb",x"49"),
   330 => (x"98",x"70",x"86",x"c4"),
   331 => (x"c0",x"87",x"c5",x"05"),
   332 => (x"87",x"ce",x"c9",x"48"),
   333 => (x"7e",x"c1",x"4d",x"c0"),
   334 => (x"bf",x"db",x"f2",x"c0"),
   335 => (x"ec",x"e3",x"c2",x"49"),
   336 => (x"4b",x"c8",x"71",x"4a"),
   337 => (x"70",x"87",x"fd",x"ec"),
   338 => (x"87",x"c2",x"05",x"98"),
   339 => (x"f2",x"c0",x"7e",x"c0"),
   340 => (x"c2",x"49",x"bf",x"d7"),
   341 => (x"71",x"4a",x"c8",x"e4"),
   342 => (x"e7",x"ec",x"4b",x"c8"),
   343 => (x"05",x"98",x"70",x"87"),
   344 => (x"7e",x"c0",x"87",x"c2"),
   345 => (x"fd",x"c0",x"02",x"6e"),
   346 => (x"fc",x"e9",x"c2",x"87"),
   347 => (x"ea",x"c2",x"4d",x"bf"),
   348 => (x"7e",x"bf",x"9f",x"f4"),
   349 => (x"ea",x"d6",x"c5",x"48"),
   350 => (x"87",x"c7",x"05",x"a8"),
   351 => (x"bf",x"fc",x"e9",x"c2"),
   352 => (x"6e",x"87",x"ce",x"4d"),
   353 => (x"d5",x"e9",x"ca",x"48"),
   354 => (x"87",x"c5",x"02",x"a8"),
   355 => (x"f1",x"c7",x"48",x"c0"),
   356 => (x"f6",x"e2",x"c2",x"87"),
   357 => (x"f9",x"49",x"75",x"1e"),
   358 => (x"86",x"c4",x"87",x"ec"),
   359 => (x"c5",x"05",x"98",x"70"),
   360 => (x"c7",x"48",x"c0",x"87"),
   361 => (x"f2",x"c0",x"87",x"dc"),
   362 => (x"c2",x"49",x"bf",x"d7"),
   363 => (x"71",x"4a",x"c8",x"e4"),
   364 => (x"cf",x"eb",x"4b",x"c8"),
   365 => (x"05",x"98",x"70",x"87"),
   366 => (x"ea",x"c2",x"87",x"c8"),
   367 => (x"78",x"c1",x"48",x"fe"),
   368 => (x"f2",x"c0",x"87",x"da"),
   369 => (x"c2",x"49",x"bf",x"db"),
   370 => (x"71",x"4a",x"ec",x"e3"),
   371 => (x"f3",x"ea",x"4b",x"c8"),
   372 => (x"02",x"98",x"70",x"87"),
   373 => (x"c0",x"87",x"c5",x"c0"),
   374 => (x"87",x"e6",x"c6",x"48"),
   375 => (x"97",x"f4",x"ea",x"c2"),
   376 => (x"d5",x"c1",x"49",x"bf"),
   377 => (x"cd",x"c0",x"05",x"a9"),
   378 => (x"f5",x"ea",x"c2",x"87"),
   379 => (x"c2",x"49",x"bf",x"97"),
   380 => (x"c0",x"02",x"a9",x"ea"),
   381 => (x"48",x"c0",x"87",x"c5"),
   382 => (x"c2",x"87",x"c7",x"c6"),
   383 => (x"bf",x"97",x"f6",x"e2"),
   384 => (x"e9",x"c3",x"48",x"7e"),
   385 => (x"ce",x"c0",x"02",x"a8"),
   386 => (x"c3",x"48",x"6e",x"87"),
   387 => (x"c0",x"02",x"a8",x"eb"),
   388 => (x"48",x"c0",x"87",x"c5"),
   389 => (x"c2",x"87",x"eb",x"c5"),
   390 => (x"bf",x"97",x"c1",x"e3"),
   391 => (x"c0",x"05",x"99",x"49"),
   392 => (x"e3",x"c2",x"87",x"cc"),
   393 => (x"49",x"bf",x"97",x"c2"),
   394 => (x"c0",x"02",x"a9",x"c2"),
   395 => (x"48",x"c0",x"87",x"c5"),
   396 => (x"c2",x"87",x"cf",x"c5"),
   397 => (x"bf",x"97",x"c3",x"e3"),
   398 => (x"fa",x"ea",x"c2",x"48"),
   399 => (x"48",x"4c",x"70",x"58"),
   400 => (x"ea",x"c2",x"88",x"c1"),
   401 => (x"e3",x"c2",x"58",x"fe"),
   402 => (x"49",x"bf",x"97",x"c4"),
   403 => (x"e3",x"c2",x"81",x"75"),
   404 => (x"4a",x"bf",x"97",x"c5"),
   405 => (x"a1",x"72",x"32",x"c8"),
   406 => (x"cb",x"ef",x"c2",x"7e"),
   407 => (x"c2",x"78",x"6e",x"48"),
   408 => (x"bf",x"97",x"c6",x"e3"),
   409 => (x"58",x"a6",x"c8",x"48"),
   410 => (x"bf",x"fe",x"ea",x"c2"),
   411 => (x"87",x"d4",x"c2",x"02"),
   412 => (x"bf",x"d7",x"f2",x"c0"),
   413 => (x"c8",x"e4",x"c2",x"49"),
   414 => (x"4b",x"c8",x"71",x"4a"),
   415 => (x"70",x"87",x"c5",x"e8"),
   416 => (x"c5",x"c0",x"02",x"98"),
   417 => (x"c3",x"48",x"c0",x"87"),
   418 => (x"ea",x"c2",x"87",x"f8"),
   419 => (x"c2",x"4c",x"bf",x"f6"),
   420 => (x"c2",x"5c",x"df",x"ef"),
   421 => (x"bf",x"97",x"db",x"e3"),
   422 => (x"c2",x"31",x"c8",x"49"),
   423 => (x"bf",x"97",x"da",x"e3"),
   424 => (x"c2",x"49",x"a1",x"4a"),
   425 => (x"bf",x"97",x"dc",x"e3"),
   426 => (x"72",x"32",x"d0",x"4a"),
   427 => (x"e3",x"c2",x"49",x"a1"),
   428 => (x"4a",x"bf",x"97",x"dd"),
   429 => (x"a1",x"72",x"32",x"d8"),
   430 => (x"91",x"66",x"c4",x"49"),
   431 => (x"bf",x"cb",x"ef",x"c2"),
   432 => (x"d3",x"ef",x"c2",x"81"),
   433 => (x"e3",x"e3",x"c2",x"59"),
   434 => (x"c8",x"4a",x"bf",x"97"),
   435 => (x"e2",x"e3",x"c2",x"32"),
   436 => (x"a2",x"4b",x"bf",x"97"),
   437 => (x"e4",x"e3",x"c2",x"4a"),
   438 => (x"d0",x"4b",x"bf",x"97"),
   439 => (x"4a",x"a2",x"73",x"33"),
   440 => (x"97",x"e5",x"e3",x"c2"),
   441 => (x"9b",x"cf",x"4b",x"bf"),
   442 => (x"a2",x"73",x"33",x"d8"),
   443 => (x"d7",x"ef",x"c2",x"4a"),
   444 => (x"d3",x"ef",x"c2",x"5a"),
   445 => (x"8a",x"c2",x"4a",x"bf"),
   446 => (x"ef",x"c2",x"92",x"74"),
   447 => (x"a1",x"72",x"48",x"d7"),
   448 => (x"87",x"ca",x"c1",x"78"),
   449 => (x"97",x"c8",x"e3",x"c2"),
   450 => (x"31",x"c8",x"49",x"bf"),
   451 => (x"97",x"c7",x"e3",x"c2"),
   452 => (x"49",x"a1",x"4a",x"bf"),
   453 => (x"59",x"c6",x"eb",x"c2"),
   454 => (x"bf",x"c2",x"eb",x"c2"),
   455 => (x"c7",x"31",x"c5",x"49"),
   456 => (x"29",x"c9",x"81",x"ff"),
   457 => (x"59",x"df",x"ef",x"c2"),
   458 => (x"97",x"cd",x"e3",x"c2"),
   459 => (x"32",x"c8",x"4a",x"bf"),
   460 => (x"97",x"cc",x"e3",x"c2"),
   461 => (x"4a",x"a2",x"4b",x"bf"),
   462 => (x"6e",x"92",x"66",x"c4"),
   463 => (x"db",x"ef",x"c2",x"82"),
   464 => (x"d3",x"ef",x"c2",x"5a"),
   465 => (x"c2",x"78",x"c0",x"48"),
   466 => (x"72",x"48",x"cf",x"ef"),
   467 => (x"ef",x"c2",x"78",x"a1"),
   468 => (x"ef",x"c2",x"48",x"df"),
   469 => (x"c2",x"78",x"bf",x"d3"),
   470 => (x"c2",x"48",x"e3",x"ef"),
   471 => (x"78",x"bf",x"d7",x"ef"),
   472 => (x"bf",x"fe",x"ea",x"c2"),
   473 => (x"87",x"c9",x"c0",x"02"),
   474 => (x"30",x"c4",x"48",x"74"),
   475 => (x"c9",x"c0",x"7e",x"70"),
   476 => (x"db",x"ef",x"c2",x"87"),
   477 => (x"30",x"c4",x"48",x"bf"),
   478 => (x"eb",x"c2",x"7e",x"70"),
   479 => (x"78",x"6e",x"48",x"c2"),
   480 => (x"8e",x"f8",x"48",x"c1"),
   481 => (x"4c",x"26",x"4d",x"26"),
   482 => (x"4f",x"26",x"4b",x"26"),
   483 => (x"5c",x"5b",x"5e",x"0e"),
   484 => (x"4a",x"71",x"0e",x"5d"),
   485 => (x"bf",x"fe",x"ea",x"c2"),
   486 => (x"72",x"87",x"cb",x"02"),
   487 => (x"72",x"2b",x"c7",x"4b"),
   488 => (x"9c",x"ff",x"c1",x"4c"),
   489 => (x"4b",x"72",x"87",x"c9"),
   490 => (x"4c",x"72",x"2b",x"c8"),
   491 => (x"c2",x"9c",x"ff",x"c3"),
   492 => (x"83",x"bf",x"cb",x"ef"),
   493 => (x"bf",x"d3",x"f2",x"c0"),
   494 => (x"87",x"d9",x"02",x"ab"),
   495 => (x"5b",x"d7",x"f2",x"c0"),
   496 => (x"1e",x"f6",x"e2",x"c2"),
   497 => (x"fd",x"f0",x"49",x"73"),
   498 => (x"70",x"86",x"c4",x"87"),
   499 => (x"87",x"c5",x"05",x"98"),
   500 => (x"e6",x"c0",x"48",x"c0"),
   501 => (x"fe",x"ea",x"c2",x"87"),
   502 => (x"87",x"d2",x"02",x"bf"),
   503 => (x"91",x"c4",x"49",x"74"),
   504 => (x"81",x"f6",x"e2",x"c2"),
   505 => (x"ff",x"cf",x"4d",x"69"),
   506 => (x"9d",x"ff",x"ff",x"ff"),
   507 => (x"49",x"74",x"87",x"cb"),
   508 => (x"e2",x"c2",x"91",x"c2"),
   509 => (x"69",x"9f",x"81",x"f6"),
   510 => (x"fe",x"48",x"75",x"4d"),
   511 => (x"5e",x"0e",x"87",x"c6"),
   512 => (x"0e",x"5d",x"5c",x"5b"),
   513 => (x"c0",x"4d",x"71",x"1e"),
   514 => (x"ca",x"49",x"c1",x"1e"),
   515 => (x"86",x"c4",x"87",x"ee"),
   516 => (x"02",x"9c",x"4c",x"70"),
   517 => (x"c2",x"87",x"c0",x"c1"),
   518 => (x"75",x"4a",x"c6",x"eb"),
   519 => (x"87",x"c9",x"e1",x"49"),
   520 => (x"c0",x"02",x"98",x"70"),
   521 => (x"4a",x"74",x"87",x"f1"),
   522 => (x"4b",x"cb",x"49",x"75"),
   523 => (x"70",x"87",x"ef",x"e1"),
   524 => (x"e2",x"c0",x"02",x"98"),
   525 => (x"74",x"1e",x"c0",x"87"),
   526 => (x"87",x"c7",x"02",x"9c"),
   527 => (x"c0",x"48",x"a6",x"c4"),
   528 => (x"c4",x"87",x"c5",x"78"),
   529 => (x"78",x"c1",x"48",x"a6"),
   530 => (x"c9",x"49",x"66",x"c4"),
   531 => (x"86",x"c4",x"87",x"ee"),
   532 => (x"05",x"9c",x"4c",x"70"),
   533 => (x"74",x"87",x"c0",x"ff"),
   534 => (x"e7",x"fc",x"26",x"48"),
   535 => (x"5b",x"5e",x"0e",x"87"),
   536 => (x"1e",x"0e",x"5d",x"5c"),
   537 => (x"05",x"9b",x"4b",x"71"),
   538 => (x"48",x"c0",x"87",x"c5"),
   539 => (x"c8",x"87",x"e5",x"c1"),
   540 => (x"7d",x"c0",x"4d",x"a3"),
   541 => (x"c7",x"02",x"66",x"d4"),
   542 => (x"97",x"66",x"d4",x"87"),
   543 => (x"87",x"c5",x"05",x"bf"),
   544 => (x"cf",x"c1",x"48",x"c0"),
   545 => (x"49",x"66",x"d4",x"87"),
   546 => (x"70",x"87",x"f3",x"fd"),
   547 => (x"c1",x"02",x"9c",x"4c"),
   548 => (x"a4",x"dc",x"87",x"c0"),
   549 => (x"da",x"7d",x"69",x"49"),
   550 => (x"a3",x"c4",x"49",x"a4"),
   551 => (x"7a",x"69",x"9f",x"4a"),
   552 => (x"bf",x"fe",x"ea",x"c2"),
   553 => (x"d4",x"87",x"d2",x"02"),
   554 => (x"69",x"9f",x"49",x"a4"),
   555 => (x"ff",x"ff",x"c0",x"49"),
   556 => (x"d0",x"48",x"71",x"99"),
   557 => (x"c2",x"7e",x"70",x"30"),
   558 => (x"6e",x"7e",x"c0",x"87"),
   559 => (x"80",x"6a",x"48",x"49"),
   560 => (x"7b",x"c0",x"7a",x"70"),
   561 => (x"6a",x"49",x"a3",x"cc"),
   562 => (x"49",x"a3",x"d0",x"79"),
   563 => (x"48",x"74",x"79",x"c0"),
   564 => (x"48",x"c0",x"87",x"c2"),
   565 => (x"87",x"ec",x"fa",x"26"),
   566 => (x"5c",x"5b",x"5e",x"0e"),
   567 => (x"4c",x"71",x"0e",x"5d"),
   568 => (x"48",x"d3",x"f2",x"c0"),
   569 => (x"9c",x"74",x"78",x"ff"),
   570 => (x"87",x"ca",x"c1",x"02"),
   571 => (x"69",x"49",x"a4",x"c8"),
   572 => (x"87",x"c2",x"c1",x"02"),
   573 => (x"6c",x"4a",x"66",x"d0"),
   574 => (x"a6",x"d4",x"82",x"49"),
   575 => (x"4d",x"66",x"d0",x"5a"),
   576 => (x"fa",x"ea",x"c2",x"b9"),
   577 => (x"ba",x"ff",x"4a",x"bf"),
   578 => (x"99",x"71",x"99",x"72"),
   579 => (x"87",x"e4",x"c0",x"02"),
   580 => (x"6b",x"4b",x"a4",x"c4"),
   581 => (x"87",x"f4",x"f9",x"49"),
   582 => (x"ea",x"c2",x"7b",x"70"),
   583 => (x"6c",x"49",x"bf",x"f6"),
   584 => (x"75",x"7c",x"71",x"81"),
   585 => (x"fa",x"ea",x"c2",x"b9"),
   586 => (x"ba",x"ff",x"4a",x"bf"),
   587 => (x"99",x"71",x"99",x"72"),
   588 => (x"87",x"dc",x"ff",x"05"),
   589 => (x"cb",x"f9",x"7c",x"75"),
   590 => (x"1e",x"73",x"1e",x"87"),
   591 => (x"02",x"9b",x"4b",x"71"),
   592 => (x"a3",x"c8",x"87",x"c7"),
   593 => (x"c5",x"05",x"69",x"49"),
   594 => (x"c0",x"48",x"c0",x"87"),
   595 => (x"ef",x"c2",x"87",x"eb"),
   596 => (x"c4",x"4a",x"bf",x"cf"),
   597 => (x"49",x"69",x"49",x"a3"),
   598 => (x"ea",x"c2",x"89",x"c2"),
   599 => (x"71",x"91",x"bf",x"f6"),
   600 => (x"ea",x"c2",x"4a",x"a2"),
   601 => (x"6b",x"49",x"bf",x"fa"),
   602 => (x"4a",x"a2",x"71",x"99"),
   603 => (x"72",x"1e",x"66",x"c8"),
   604 => (x"87",x"d2",x"ea",x"49"),
   605 => (x"49",x"70",x"86",x"c4"),
   606 => (x"87",x"cc",x"f8",x"48"),
   607 => (x"71",x"1e",x"73",x"1e"),
   608 => (x"c7",x"02",x"9b",x"4b"),
   609 => (x"49",x"a3",x"c8",x"87"),
   610 => (x"87",x"c5",x"05",x"69"),
   611 => (x"eb",x"c0",x"48",x"c0"),
   612 => (x"cf",x"ef",x"c2",x"87"),
   613 => (x"a3",x"c4",x"4a",x"bf"),
   614 => (x"c2",x"49",x"69",x"49"),
   615 => (x"f6",x"ea",x"c2",x"89"),
   616 => (x"a2",x"71",x"91",x"bf"),
   617 => (x"fa",x"ea",x"c2",x"4a"),
   618 => (x"99",x"6b",x"49",x"bf"),
   619 => (x"c8",x"4a",x"a2",x"71"),
   620 => (x"49",x"72",x"1e",x"66"),
   621 => (x"c4",x"87",x"c5",x"e6"),
   622 => (x"48",x"49",x"70",x"86"),
   623 => (x"0e",x"87",x"c9",x"f7"),
   624 => (x"5d",x"5c",x"5b",x"5e"),
   625 => (x"4b",x"71",x"1e",x"0e"),
   626 => (x"c9",x"4c",x"66",x"d4"),
   627 => (x"02",x"9b",x"73",x"2c"),
   628 => (x"c8",x"87",x"cf",x"c1"),
   629 => (x"02",x"69",x"49",x"a3"),
   630 => (x"d0",x"87",x"c7",x"c1"),
   631 => (x"66",x"d4",x"4d",x"a3"),
   632 => (x"fa",x"ea",x"c2",x"7d"),
   633 => (x"b9",x"ff",x"49",x"bf"),
   634 => (x"7e",x"99",x"4a",x"6b"),
   635 => (x"cd",x"03",x"ac",x"71"),
   636 => (x"7d",x"7b",x"c0",x"87"),
   637 => (x"c4",x"4a",x"a3",x"cc"),
   638 => (x"79",x"6a",x"49",x"a3"),
   639 => (x"8c",x"72",x"87",x"c2"),
   640 => (x"dd",x"02",x"9c",x"74"),
   641 => (x"73",x"1e",x"49",x"87"),
   642 => (x"87",x"cc",x"fb",x"49"),
   643 => (x"66",x"d4",x"86",x"c4"),
   644 => (x"99",x"ff",x"c7",x"49"),
   645 => (x"c2",x"87",x"cb",x"02"),
   646 => (x"73",x"1e",x"f6",x"e2"),
   647 => (x"87",x"d9",x"fc",x"49"),
   648 => (x"f5",x"26",x"86",x"c4"),
   649 => (x"73",x"1e",x"87",x"de"),
   650 => (x"9b",x"4b",x"71",x"1e"),
   651 => (x"87",x"e4",x"c0",x"02"),
   652 => (x"5b",x"e3",x"ef",x"c2"),
   653 => (x"8a",x"c2",x"4a",x"73"),
   654 => (x"bf",x"f6",x"ea",x"c2"),
   655 => (x"ef",x"c2",x"92",x"49"),
   656 => (x"72",x"48",x"bf",x"cf"),
   657 => (x"e7",x"ef",x"c2",x"80"),
   658 => (x"c4",x"48",x"71",x"58"),
   659 => (x"c6",x"eb",x"c2",x"30"),
   660 => (x"87",x"ed",x"c0",x"58"),
   661 => (x"48",x"df",x"ef",x"c2"),
   662 => (x"bf",x"d3",x"ef",x"c2"),
   663 => (x"e3",x"ef",x"c2",x"78"),
   664 => (x"d7",x"ef",x"c2",x"48"),
   665 => (x"ea",x"c2",x"78",x"bf"),
   666 => (x"c9",x"02",x"bf",x"fe"),
   667 => (x"f6",x"ea",x"c2",x"87"),
   668 => (x"31",x"c4",x"49",x"bf"),
   669 => (x"ef",x"c2",x"87",x"c7"),
   670 => (x"c4",x"49",x"bf",x"db"),
   671 => (x"c6",x"eb",x"c2",x"31"),
   672 => (x"87",x"c4",x"f4",x"59"),
   673 => (x"5c",x"5b",x"5e",x"0e"),
   674 => (x"c0",x"4a",x"71",x"0e"),
   675 => (x"02",x"9a",x"72",x"4b"),
   676 => (x"da",x"87",x"e1",x"c0"),
   677 => (x"69",x"9f",x"49",x"a2"),
   678 => (x"fe",x"ea",x"c2",x"4b"),
   679 => (x"87",x"cf",x"02",x"bf"),
   680 => (x"9f",x"49",x"a2",x"d4"),
   681 => (x"c0",x"4c",x"49",x"69"),
   682 => (x"d0",x"9c",x"ff",x"ff"),
   683 => (x"c0",x"87",x"c2",x"34"),
   684 => (x"b3",x"49",x"74",x"4c"),
   685 => (x"ed",x"fd",x"49",x"73"),
   686 => (x"87",x"ca",x"f3",x"87"),
   687 => (x"5c",x"5b",x"5e",x"0e"),
   688 => (x"86",x"f4",x"0e",x"5d"),
   689 => (x"7e",x"c0",x"4a",x"71"),
   690 => (x"d8",x"02",x"9a",x"72"),
   691 => (x"f2",x"e2",x"c2",x"87"),
   692 => (x"c2",x"78",x"c0",x"48"),
   693 => (x"c2",x"48",x"ea",x"e2"),
   694 => (x"78",x"bf",x"e3",x"ef"),
   695 => (x"48",x"ee",x"e2",x"c2"),
   696 => (x"bf",x"df",x"ef",x"c2"),
   697 => (x"d3",x"eb",x"c2",x"78"),
   698 => (x"c2",x"50",x"c0",x"48"),
   699 => (x"49",x"bf",x"c2",x"eb"),
   700 => (x"bf",x"f2",x"e2",x"c2"),
   701 => (x"03",x"aa",x"71",x"4a"),
   702 => (x"72",x"87",x"ff",x"c3"),
   703 => (x"05",x"99",x"cf",x"49"),
   704 => (x"c2",x"87",x"e0",x"c0"),
   705 => (x"c2",x"1e",x"f6",x"e2"),
   706 => (x"49",x"bf",x"ea",x"e2"),
   707 => (x"48",x"ea",x"e2",x"c2"),
   708 => (x"71",x"78",x"a1",x"c1"),
   709 => (x"c4",x"87",x"ef",x"e3"),
   710 => (x"cf",x"f2",x"c0",x"86"),
   711 => (x"f6",x"e2",x"c2",x"48"),
   712 => (x"c0",x"87",x"cc",x"78"),
   713 => (x"48",x"bf",x"cf",x"f2"),
   714 => (x"c0",x"80",x"e0",x"c0"),
   715 => (x"c2",x"58",x"d3",x"f2"),
   716 => (x"48",x"bf",x"f2",x"e2"),
   717 => (x"e2",x"c2",x"80",x"c1"),
   718 => (x"8f",x"27",x"58",x"f6"),
   719 => (x"bf",x"00",x"00",x"0c"),
   720 => (x"9d",x"4d",x"bf",x"97"),
   721 => (x"87",x"e2",x"c2",x"02"),
   722 => (x"02",x"ad",x"e5",x"c3"),
   723 => (x"c0",x"87",x"db",x"c2"),
   724 => (x"4b",x"bf",x"cf",x"f2"),
   725 => (x"11",x"49",x"a3",x"cb"),
   726 => (x"05",x"ac",x"cf",x"4c"),
   727 => (x"75",x"87",x"d2",x"c1"),
   728 => (x"c1",x"99",x"df",x"49"),
   729 => (x"c2",x"91",x"cd",x"89"),
   730 => (x"c1",x"81",x"c6",x"eb"),
   731 => (x"51",x"12",x"4a",x"a3"),
   732 => (x"12",x"4a",x"a3",x"c3"),
   733 => (x"4a",x"a3",x"c5",x"51"),
   734 => (x"a3",x"c7",x"51",x"12"),
   735 => (x"c9",x"51",x"12",x"4a"),
   736 => (x"51",x"12",x"4a",x"a3"),
   737 => (x"12",x"4a",x"a3",x"ce"),
   738 => (x"4a",x"a3",x"d0",x"51"),
   739 => (x"a3",x"d2",x"51",x"12"),
   740 => (x"d4",x"51",x"12",x"4a"),
   741 => (x"51",x"12",x"4a",x"a3"),
   742 => (x"12",x"4a",x"a3",x"d6"),
   743 => (x"4a",x"a3",x"d8",x"51"),
   744 => (x"a3",x"dc",x"51",x"12"),
   745 => (x"de",x"51",x"12",x"4a"),
   746 => (x"51",x"12",x"4a",x"a3"),
   747 => (x"f9",x"c0",x"7e",x"c1"),
   748 => (x"c8",x"49",x"74",x"87"),
   749 => (x"ea",x"c0",x"05",x"99"),
   750 => (x"d0",x"49",x"74",x"87"),
   751 => (x"87",x"d0",x"05",x"99"),
   752 => (x"c0",x"02",x"66",x"dc"),
   753 => (x"49",x"73",x"87",x"ca"),
   754 => (x"70",x"0f",x"66",x"dc"),
   755 => (x"87",x"d3",x"02",x"98"),
   756 => (x"c6",x"c0",x"05",x"6e"),
   757 => (x"c6",x"eb",x"c2",x"87"),
   758 => (x"c0",x"50",x"c0",x"48"),
   759 => (x"48",x"bf",x"cf",x"f2"),
   760 => (x"c2",x"87",x"e7",x"c2"),
   761 => (x"c0",x"48",x"d3",x"eb"),
   762 => (x"eb",x"c2",x"7e",x"50"),
   763 => (x"c2",x"49",x"bf",x"c2"),
   764 => (x"4a",x"bf",x"f2",x"e2"),
   765 => (x"fc",x"04",x"aa",x"71"),
   766 => (x"ef",x"c2",x"87",x"c1"),
   767 => (x"c0",x"05",x"bf",x"e3"),
   768 => (x"ea",x"c2",x"87",x"c8"),
   769 => (x"c1",x"02",x"bf",x"fe"),
   770 => (x"f2",x"c0",x"87",x"fe"),
   771 => (x"78",x"ff",x"48",x"d3"),
   772 => (x"bf",x"ee",x"e2",x"c2"),
   773 => (x"87",x"f4",x"ed",x"49"),
   774 => (x"e2",x"c2",x"49",x"70"),
   775 => (x"a6",x"c4",x"59",x"f2"),
   776 => (x"ee",x"e2",x"c2",x"48"),
   777 => (x"ea",x"c2",x"78",x"bf"),
   778 => (x"c0",x"02",x"bf",x"fe"),
   779 => (x"66",x"c4",x"87",x"d8"),
   780 => (x"ff",x"ff",x"cf",x"49"),
   781 => (x"a9",x"99",x"f8",x"ff"),
   782 => (x"87",x"c5",x"c0",x"02"),
   783 => (x"e1",x"c0",x"4d",x"c0"),
   784 => (x"c0",x"4d",x"c1",x"87"),
   785 => (x"66",x"c4",x"87",x"dc"),
   786 => (x"f8",x"ff",x"cf",x"49"),
   787 => (x"c0",x"02",x"a9",x"99"),
   788 => (x"a6",x"c8",x"87",x"c8"),
   789 => (x"c0",x"78",x"c0",x"48"),
   790 => (x"a6",x"c8",x"87",x"c5"),
   791 => (x"c8",x"78",x"c1",x"48"),
   792 => (x"9d",x"75",x"4d",x"66"),
   793 => (x"87",x"e0",x"c0",x"05"),
   794 => (x"c2",x"49",x"66",x"c4"),
   795 => (x"f6",x"ea",x"c2",x"89"),
   796 => (x"c2",x"91",x"4a",x"bf"),
   797 => (x"4a",x"bf",x"cf",x"ef"),
   798 => (x"48",x"ea",x"e2",x"c2"),
   799 => (x"c2",x"78",x"a1",x"72"),
   800 => (x"c0",x"48",x"f2",x"e2"),
   801 => (x"87",x"e3",x"f9",x"78"),
   802 => (x"8e",x"f4",x"48",x"c0"),
   803 => (x"00",x"87",x"f5",x"eb"),
   804 => (x"ff",x"00",x"00",x"00"),
   805 => (x"9f",x"ff",x"ff",x"ff"),
   806 => (x"a8",x"00",x"00",x"0c"),
   807 => (x"46",x"00",x"00",x"0c"),
   808 => (x"32",x"33",x"54",x"41"),
   809 => (x"00",x"20",x"20",x"20"),
   810 => (x"31",x"54",x"41",x"46"),
   811 => (x"20",x"20",x"20",x"36"),
   812 => (x"d4",x"ff",x"1e",x"00"),
   813 => (x"78",x"ff",x"c3",x"48"),
   814 => (x"4f",x"26",x"48",x"68"),
   815 => (x"48",x"d4",x"ff",x"1e"),
   816 => (x"ff",x"78",x"ff",x"c3"),
   817 => (x"e1",x"c8",x"48",x"d0"),
   818 => (x"48",x"d4",x"ff",x"78"),
   819 => (x"ef",x"c2",x"78",x"d4"),
   820 => (x"d4",x"ff",x"48",x"e7"),
   821 => (x"4f",x"26",x"50",x"bf"),
   822 => (x"48",x"d0",x"ff",x"1e"),
   823 => (x"26",x"78",x"e0",x"c0"),
   824 => (x"cc",x"ff",x"1e",x"4f"),
   825 => (x"99",x"49",x"70",x"87"),
   826 => (x"c0",x"87",x"c6",x"02"),
   827 => (x"f1",x"05",x"a9",x"fb"),
   828 => (x"26",x"48",x"71",x"87"),
   829 => (x"5b",x"5e",x"0e",x"4f"),
   830 => (x"4b",x"71",x"0e",x"5c"),
   831 => (x"f0",x"fe",x"4c",x"c0"),
   832 => (x"99",x"49",x"70",x"87"),
   833 => (x"87",x"f9",x"c0",x"02"),
   834 => (x"02",x"a9",x"ec",x"c0"),
   835 => (x"c0",x"87",x"f2",x"c0"),
   836 => (x"c0",x"02",x"a9",x"fb"),
   837 => (x"66",x"cc",x"87",x"eb"),
   838 => (x"c7",x"03",x"ac",x"b7"),
   839 => (x"02",x"66",x"d0",x"87"),
   840 => (x"53",x"71",x"87",x"c2"),
   841 => (x"c2",x"02",x"99",x"71"),
   842 => (x"fe",x"84",x"c1",x"87"),
   843 => (x"49",x"70",x"87",x"c3"),
   844 => (x"87",x"cd",x"02",x"99"),
   845 => (x"02",x"a9",x"ec",x"c0"),
   846 => (x"fb",x"c0",x"87",x"c7"),
   847 => (x"d5",x"ff",x"05",x"a9"),
   848 => (x"02",x"66",x"d0",x"87"),
   849 => (x"97",x"c0",x"87",x"c3"),
   850 => (x"a9",x"ec",x"c0",x"7b"),
   851 => (x"74",x"87",x"c4",x"05"),
   852 => (x"74",x"87",x"c5",x"4a"),
   853 => (x"8a",x"0a",x"c0",x"4a"),
   854 => (x"87",x"c2",x"48",x"72"),
   855 => (x"4c",x"26",x"4d",x"26"),
   856 => (x"4f",x"26",x"4b",x"26"),
   857 => (x"87",x"c9",x"fd",x"1e"),
   858 => (x"f0",x"c0",x"49",x"70"),
   859 => (x"ca",x"04",x"a9",x"b7"),
   860 => (x"b7",x"f9",x"c0",x"87"),
   861 => (x"87",x"c3",x"01",x"a9"),
   862 => (x"c1",x"89",x"f0",x"c0"),
   863 => (x"04",x"a9",x"b7",x"c1"),
   864 => (x"da",x"c1",x"87",x"ca"),
   865 => (x"c3",x"01",x"a9",x"b7"),
   866 => (x"89",x"f7",x"c0",x"87"),
   867 => (x"4f",x"26",x"48",x"71"),
   868 => (x"5c",x"5b",x"5e",x"0e"),
   869 => (x"ff",x"4a",x"71",x"0e"),
   870 => (x"49",x"72",x"4c",x"d4"),
   871 => (x"70",x"87",x"ea",x"c0"),
   872 => (x"c2",x"02",x"9b",x"4b"),
   873 => (x"ff",x"8b",x"c1",x"87"),
   874 => (x"c5",x"c8",x"48",x"d0"),
   875 => (x"7c",x"d5",x"c1",x"78"),
   876 => (x"31",x"c6",x"49",x"73"),
   877 => (x"97",x"ec",x"de",x"c2"),
   878 => (x"71",x"48",x"4a",x"bf"),
   879 => (x"ff",x"7c",x"70",x"b0"),
   880 => (x"78",x"c4",x"48",x"d0"),
   881 => (x"d5",x"fe",x"48",x"73"),
   882 => (x"5b",x"5e",x"0e",x"87"),
   883 => (x"f8",x"0e",x"5d",x"5c"),
   884 => (x"c0",x"4b",x"71",x"86"),
   885 => (x"f0",x"fa",x"c0",x"7e"),
   886 => (x"df",x"49",x"bf",x"97"),
   887 => (x"ee",x"c0",x"05",x"a9"),
   888 => (x"49",x"a3",x"c8",x"87"),
   889 => (x"c1",x"49",x"69",x"97"),
   890 => (x"dd",x"05",x"a9",x"c3"),
   891 => (x"49",x"a3",x"c9",x"87"),
   892 => (x"c1",x"49",x"69",x"97"),
   893 => (x"d1",x"05",x"a9",x"c6"),
   894 => (x"49",x"a3",x"ca",x"87"),
   895 => (x"c1",x"49",x"69",x"97"),
   896 => (x"c5",x"05",x"a9",x"c7"),
   897 => (x"c2",x"48",x"c1",x"87"),
   898 => (x"48",x"c0",x"87",x"e1"),
   899 => (x"fa",x"87",x"dc",x"c2"),
   900 => (x"4c",x"c0",x"87",x"ea"),
   901 => (x"97",x"f0",x"fa",x"c0"),
   902 => (x"a9",x"c0",x"49",x"bf"),
   903 => (x"fa",x"87",x"cf",x"04"),
   904 => (x"84",x"c1",x"87",x"ff"),
   905 => (x"97",x"f0",x"fa",x"c0"),
   906 => (x"06",x"ac",x"49",x"bf"),
   907 => (x"fa",x"c0",x"87",x"f1"),
   908 => (x"02",x"bf",x"97",x"f0"),
   909 => (x"f8",x"f9",x"87",x"cf"),
   910 => (x"99",x"49",x"70",x"87"),
   911 => (x"c0",x"87",x"c6",x"02"),
   912 => (x"f1",x"05",x"a9",x"ec"),
   913 => (x"f9",x"4c",x"c0",x"87"),
   914 => (x"4d",x"70",x"87",x"e7"),
   915 => (x"c8",x"87",x"e2",x"f9"),
   916 => (x"dc",x"f9",x"58",x"a6"),
   917 => (x"c1",x"4a",x"70",x"87"),
   918 => (x"49",x"a3",x"c8",x"84"),
   919 => (x"ad",x"49",x"69",x"97"),
   920 => (x"c0",x"87",x"c7",x"02"),
   921 => (x"c0",x"05",x"ad",x"ff"),
   922 => (x"a3",x"c9",x"87",x"e7"),
   923 => (x"49",x"69",x"97",x"49"),
   924 => (x"02",x"a9",x"66",x"c4"),
   925 => (x"c0",x"48",x"87",x"c7"),
   926 => (x"d4",x"05",x"a8",x"ff"),
   927 => (x"49",x"a3",x"ca",x"87"),
   928 => (x"aa",x"49",x"69",x"97"),
   929 => (x"c0",x"87",x"c6",x"02"),
   930 => (x"c4",x"05",x"aa",x"ff"),
   931 => (x"d0",x"7e",x"c1",x"87"),
   932 => (x"ad",x"ec",x"c0",x"87"),
   933 => (x"c0",x"87",x"c6",x"02"),
   934 => (x"c4",x"05",x"ad",x"fb"),
   935 => (x"c1",x"4c",x"c0",x"87"),
   936 => (x"fe",x"02",x"6e",x"7e"),
   937 => (x"ef",x"f8",x"87",x"e1"),
   938 => (x"f8",x"48",x"74",x"87"),
   939 => (x"87",x"ec",x"fa",x"8e"),
   940 => (x"5b",x"5e",x"0e",x"00"),
   941 => (x"1e",x"0e",x"5d",x"5c"),
   942 => (x"4c",x"c0",x"4b",x"71"),
   943 => (x"c0",x"04",x"ab",x"4d"),
   944 => (x"f7",x"c0",x"87",x"e8"),
   945 => (x"9d",x"75",x"1e",x"c9"),
   946 => (x"c0",x"87",x"c4",x"02"),
   947 => (x"c1",x"87",x"c2",x"4a"),
   948 => (x"ef",x"49",x"72",x"4a"),
   949 => (x"86",x"c4",x"87",x"e6"),
   950 => (x"84",x"c1",x"7e",x"70"),
   951 => (x"87",x"c2",x"05",x"6e"),
   952 => (x"85",x"c1",x"4c",x"73"),
   953 => (x"ff",x"06",x"ac",x"73"),
   954 => (x"48",x"6e",x"87",x"d8"),
   955 => (x"26",x"4d",x"26",x"26"),
   956 => (x"26",x"4b",x"26",x"4c"),
   957 => (x"5b",x"5e",x"0e",x"4f"),
   958 => (x"1e",x"0e",x"5d",x"5c"),
   959 => (x"de",x"49",x"4c",x"71"),
   960 => (x"c1",x"f0",x"c2",x"91"),
   961 => (x"97",x"85",x"71",x"4d"),
   962 => (x"dd",x"c1",x"02",x"6d"),
   963 => (x"ec",x"ef",x"c2",x"87"),
   964 => (x"82",x"74",x"4a",x"bf"),
   965 => (x"d8",x"fe",x"49",x"72"),
   966 => (x"6e",x"7e",x"70",x"87"),
   967 => (x"87",x"f3",x"c0",x"02"),
   968 => (x"4b",x"f4",x"ef",x"c2"),
   969 => (x"49",x"cb",x"4a",x"6e"),
   970 => (x"87",x"d6",x"c6",x"ff"),
   971 => (x"93",x"cb",x"4b",x"74"),
   972 => (x"83",x"e0",x"e1",x"c1"),
   973 => (x"fd",x"c0",x"83",x"c4"),
   974 => (x"49",x"74",x"7b",x"ee"),
   975 => (x"87",x"f7",x"c5",x"c1"),
   976 => (x"f0",x"c2",x"7b",x"75"),
   977 => (x"49",x"bf",x"97",x"c0"),
   978 => (x"f4",x"ef",x"c2",x"1e"),
   979 => (x"f9",x"df",x"c1",x"49"),
   980 => (x"74",x"86",x"c4",x"87"),
   981 => (x"de",x"c5",x"c1",x"49"),
   982 => (x"c1",x"49",x"c0",x"87"),
   983 => (x"c2",x"87",x"fd",x"c6"),
   984 => (x"c0",x"48",x"e8",x"ef"),
   985 => (x"df",x"49",x"c1",x"78"),
   986 => (x"fd",x"26",x"87",x"fd"),
   987 => (x"6f",x"4c",x"87",x"ff"),
   988 => (x"6e",x"69",x"64",x"61"),
   989 => (x"2e",x"2e",x"2e",x"67"),
   990 => (x"5b",x"5e",x"0e",x"00"),
   991 => (x"4b",x"71",x"0e",x"5c"),
   992 => (x"ec",x"ef",x"c2",x"4a"),
   993 => (x"49",x"72",x"82",x"bf"),
   994 => (x"70",x"87",x"e6",x"fc"),
   995 => (x"c4",x"02",x"9c",x"4c"),
   996 => (x"ef",x"eb",x"49",x"87"),
   997 => (x"ec",x"ef",x"c2",x"87"),
   998 => (x"c1",x"78",x"c0",x"48"),
   999 => (x"87",x"c7",x"df",x"49"),
  1000 => (x"0e",x"87",x"cc",x"fd"),
  1001 => (x"5d",x"5c",x"5b",x"5e"),
  1002 => (x"c2",x"86",x"f4",x"0e"),
  1003 => (x"c0",x"4d",x"f6",x"e2"),
  1004 => (x"48",x"a6",x"c4",x"4c"),
  1005 => (x"ef",x"c2",x"78",x"c0"),
  1006 => (x"c0",x"49",x"bf",x"ec"),
  1007 => (x"c1",x"c1",x"06",x"a9"),
  1008 => (x"f6",x"e2",x"c2",x"87"),
  1009 => (x"c0",x"02",x"98",x"48"),
  1010 => (x"f7",x"c0",x"87",x"f8"),
  1011 => (x"66",x"c8",x"1e",x"c9"),
  1012 => (x"c4",x"87",x"c7",x"02"),
  1013 => (x"78",x"c0",x"48",x"a6"),
  1014 => (x"a6",x"c4",x"87",x"c5"),
  1015 => (x"c4",x"78",x"c1",x"48"),
  1016 => (x"d7",x"eb",x"49",x"66"),
  1017 => (x"70",x"86",x"c4",x"87"),
  1018 => (x"c4",x"84",x"c1",x"4d"),
  1019 => (x"80",x"c1",x"48",x"66"),
  1020 => (x"c2",x"58",x"a6",x"c8"),
  1021 => (x"49",x"bf",x"ec",x"ef"),
  1022 => (x"87",x"c6",x"03",x"ac"),
  1023 => (x"ff",x"05",x"9d",x"75"),
  1024 => (x"4c",x"c0",x"87",x"c8"),
  1025 => (x"c3",x"02",x"9d",x"75"),
  1026 => (x"f7",x"c0",x"87",x"e0"),
  1027 => (x"66",x"c8",x"1e",x"c9"),
  1028 => (x"cc",x"87",x"c7",x"02"),
  1029 => (x"78",x"c0",x"48",x"a6"),
  1030 => (x"a6",x"cc",x"87",x"c5"),
  1031 => (x"cc",x"78",x"c1",x"48"),
  1032 => (x"d7",x"ea",x"49",x"66"),
  1033 => (x"70",x"86",x"c4",x"87"),
  1034 => (x"c2",x"02",x"6e",x"7e"),
  1035 => (x"49",x"6e",x"87",x"e9"),
  1036 => (x"69",x"97",x"81",x"cb"),
  1037 => (x"02",x"99",x"d0",x"49"),
  1038 => (x"c0",x"87",x"d6",x"c1"),
  1039 => (x"74",x"4a",x"f9",x"fd"),
  1040 => (x"c1",x"91",x"cb",x"49"),
  1041 => (x"72",x"81",x"e0",x"e1"),
  1042 => (x"c3",x"81",x"c8",x"79"),
  1043 => (x"49",x"74",x"51",x"ff"),
  1044 => (x"f0",x"c2",x"91",x"de"),
  1045 => (x"85",x"71",x"4d",x"c1"),
  1046 => (x"7d",x"97",x"c1",x"c2"),
  1047 => (x"c0",x"49",x"a5",x"c1"),
  1048 => (x"eb",x"c2",x"51",x"e0"),
  1049 => (x"02",x"bf",x"97",x"c6"),
  1050 => (x"84",x"c1",x"87",x"d2"),
  1051 => (x"c2",x"4b",x"a5",x"c2"),
  1052 => (x"db",x"4a",x"c6",x"eb"),
  1053 => (x"c9",x"c1",x"ff",x"49"),
  1054 => (x"87",x"db",x"c1",x"87"),
  1055 => (x"c0",x"49",x"a5",x"cd"),
  1056 => (x"c2",x"84",x"c1",x"51"),
  1057 => (x"4a",x"6e",x"4b",x"a5"),
  1058 => (x"c0",x"ff",x"49",x"cb"),
  1059 => (x"c6",x"c1",x"87",x"f4"),
  1060 => (x"f5",x"fb",x"c0",x"87"),
  1061 => (x"cb",x"49",x"74",x"4a"),
  1062 => (x"e0",x"e1",x"c1",x"91"),
  1063 => (x"c2",x"79",x"72",x"81"),
  1064 => (x"bf",x"97",x"c6",x"eb"),
  1065 => (x"74",x"87",x"d8",x"02"),
  1066 => (x"c1",x"91",x"de",x"49"),
  1067 => (x"c1",x"f0",x"c2",x"84"),
  1068 => (x"c2",x"83",x"71",x"4b"),
  1069 => (x"dd",x"4a",x"c6",x"eb"),
  1070 => (x"c5",x"c0",x"ff",x"49"),
  1071 => (x"74",x"87",x"d8",x"87"),
  1072 => (x"c2",x"93",x"de",x"4b"),
  1073 => (x"cb",x"83",x"c1",x"f0"),
  1074 => (x"51",x"c0",x"49",x"a3"),
  1075 => (x"6e",x"73",x"84",x"c1"),
  1076 => (x"fe",x"49",x"cb",x"4a"),
  1077 => (x"c4",x"87",x"eb",x"ff"),
  1078 => (x"80",x"c1",x"48",x"66"),
  1079 => (x"c7",x"58",x"a6",x"c8"),
  1080 => (x"c5",x"c0",x"03",x"ac"),
  1081 => (x"fc",x"05",x"6e",x"87"),
  1082 => (x"48",x"74",x"87",x"e0"),
  1083 => (x"fc",x"f7",x"8e",x"f4"),
  1084 => (x"1e",x"73",x"1e",x"87"),
  1085 => (x"cb",x"49",x"4b",x"71"),
  1086 => (x"e0",x"e1",x"c1",x"91"),
  1087 => (x"4a",x"a1",x"c8",x"81"),
  1088 => (x"48",x"ec",x"de",x"c2"),
  1089 => (x"a1",x"c9",x"50",x"12"),
  1090 => (x"f0",x"fa",x"c0",x"4a"),
  1091 => (x"ca",x"50",x"12",x"48"),
  1092 => (x"c0",x"f0",x"c2",x"81"),
  1093 => (x"c2",x"50",x"11",x"48"),
  1094 => (x"bf",x"97",x"c0",x"f0"),
  1095 => (x"49",x"c0",x"1e",x"49"),
  1096 => (x"87",x"e6",x"d8",x"c1"),
  1097 => (x"48",x"e8",x"ef",x"c2"),
  1098 => (x"49",x"c1",x"78",x"de"),
  1099 => (x"26",x"87",x"f8",x"d8"),
  1100 => (x"1e",x"87",x"fe",x"f6"),
  1101 => (x"cb",x"49",x"4a",x"71"),
  1102 => (x"e0",x"e1",x"c1",x"91"),
  1103 => (x"11",x"81",x"c8",x"81"),
  1104 => (x"ec",x"ef",x"c2",x"48"),
  1105 => (x"ec",x"ef",x"c2",x"58"),
  1106 => (x"c1",x"78",x"c0",x"48"),
  1107 => (x"87",x"d7",x"d8",x"49"),
  1108 => (x"c0",x"1e",x"4f",x"26"),
  1109 => (x"c3",x"ff",x"c0",x"49"),
  1110 => (x"1e",x"4f",x"26",x"87"),
  1111 => (x"d2",x"02",x"99",x"71"),
  1112 => (x"f5",x"e2",x"c1",x"87"),
  1113 => (x"f7",x"50",x"c0",x"48"),
  1114 => (x"f3",x"c4",x"c1",x"80"),
  1115 => (x"ce",x"e1",x"c1",x"40"),
  1116 => (x"c1",x"87",x"ce",x"78"),
  1117 => (x"c1",x"48",x"f1",x"e2"),
  1118 => (x"fc",x"78",x"ef",x"e0"),
  1119 => (x"d2",x"c5",x"c1",x"80"),
  1120 => (x"0e",x"4f",x"26",x"78"),
  1121 => (x"0e",x"5c",x"5b",x"5e"),
  1122 => (x"cb",x"4a",x"4c",x"71"),
  1123 => (x"e0",x"e1",x"c1",x"92"),
  1124 => (x"49",x"a2",x"c8",x"82"),
  1125 => (x"97",x"4b",x"a2",x"c9"),
  1126 => (x"97",x"1e",x"4b",x"6b"),
  1127 => (x"ca",x"1e",x"49",x"69"),
  1128 => (x"c0",x"49",x"12",x"82"),
  1129 => (x"c0",x"87",x"fe",x"e9"),
  1130 => (x"87",x"fb",x"d6",x"49"),
  1131 => (x"fc",x"c0",x"49",x"74"),
  1132 => (x"8e",x"f8",x"87",x"c5"),
  1133 => (x"1e",x"87",x"f8",x"f4"),
  1134 => (x"4b",x"71",x"1e",x"73"),
  1135 => (x"87",x"c3",x"ff",x"49"),
  1136 => (x"fe",x"fe",x"49",x"73"),
  1137 => (x"87",x"e9",x"f4",x"87"),
  1138 => (x"71",x"1e",x"73",x"1e"),
  1139 => (x"4a",x"a3",x"c6",x"4b"),
  1140 => (x"c1",x"87",x"dc",x"02"),
  1141 => (x"e4",x"c0",x"02",x"8a"),
  1142 => (x"c1",x"02",x"8a",x"87"),
  1143 => (x"02",x"8a",x"87",x"e8"),
  1144 => (x"8a",x"87",x"ca",x"c1"),
  1145 => (x"87",x"ef",x"c0",x"02"),
  1146 => (x"87",x"d9",x"02",x"8a"),
  1147 => (x"c2",x"87",x"e9",x"c1"),
  1148 => (x"df",x"48",x"e8",x"ef"),
  1149 => (x"d5",x"49",x"c1",x"78"),
  1150 => (x"e6",x"c1",x"87",x"ed"),
  1151 => (x"fc",x"49",x"c7",x"87"),
  1152 => (x"de",x"c1",x"87",x"f1"),
  1153 => (x"ec",x"ef",x"c2",x"87"),
  1154 => (x"cb",x"c1",x"02",x"bf"),
  1155 => (x"88",x"c1",x"48",x"87"),
  1156 => (x"58",x"f0",x"ef",x"c2"),
  1157 => (x"c2",x"87",x"c1",x"c1"),
  1158 => (x"02",x"bf",x"f0",x"ef"),
  1159 => (x"c2",x"87",x"f9",x"c0"),
  1160 => (x"48",x"bf",x"ec",x"ef"),
  1161 => (x"ef",x"c2",x"80",x"c1"),
  1162 => (x"eb",x"c0",x"58",x"f0"),
  1163 => (x"ec",x"ef",x"c2",x"87"),
  1164 => (x"89",x"c6",x"49",x"bf"),
  1165 => (x"59",x"f0",x"ef",x"c2"),
  1166 => (x"03",x"a9",x"b7",x"c0"),
  1167 => (x"ef",x"c2",x"87",x"da"),
  1168 => (x"78",x"c0",x"48",x"ec"),
  1169 => (x"ef",x"c2",x"87",x"d2"),
  1170 => (x"cb",x"02",x"bf",x"f0"),
  1171 => (x"ec",x"ef",x"c2",x"87"),
  1172 => (x"80",x"c6",x"48",x"bf"),
  1173 => (x"58",x"f0",x"ef",x"c2"),
  1174 => (x"ca",x"d4",x"49",x"c0"),
  1175 => (x"c0",x"49",x"73",x"87"),
  1176 => (x"f2",x"87",x"d4",x"f9"),
  1177 => (x"5e",x"0e",x"87",x"cb"),
  1178 => (x"71",x"0e",x"5c",x"5b"),
  1179 => (x"1e",x"66",x"cc",x"4c"),
  1180 => (x"93",x"cb",x"4b",x"74"),
  1181 => (x"83",x"e0",x"e1",x"c1"),
  1182 => (x"6a",x"4a",x"a3",x"c4"),
  1183 => (x"d1",x"f9",x"fe",x"49"),
  1184 => (x"f1",x"c3",x"c1",x"87"),
  1185 => (x"49",x"a3",x"c8",x"7b"),
  1186 => (x"c9",x"51",x"66",x"d4"),
  1187 => (x"66",x"d8",x"49",x"a3"),
  1188 => (x"49",x"a3",x"ca",x"51"),
  1189 => (x"26",x"51",x"66",x"dc"),
  1190 => (x"0e",x"87",x"d4",x"f1"),
  1191 => (x"5d",x"5c",x"5b",x"5e"),
  1192 => (x"86",x"d0",x"ff",x"0e"),
  1193 => (x"c8",x"59",x"a6",x"d8"),
  1194 => (x"78",x"c0",x"48",x"a6"),
  1195 => (x"c4",x"c1",x"80",x"fc"),
  1196 => (x"80",x"c8",x"78",x"66"),
  1197 => (x"80",x"c4",x"78",x"c1"),
  1198 => (x"ef",x"c2",x"78",x"c1"),
  1199 => (x"78",x"c1",x"48",x"f0"),
  1200 => (x"bf",x"e8",x"ef",x"c2"),
  1201 => (x"de",x"48",x"6e",x"7e"),
  1202 => (x"87",x"cb",x"05",x"a8"),
  1203 => (x"70",x"87",x"d4",x"f3"),
  1204 => (x"59",x"a6",x"cc",x"49"),
  1205 => (x"6e",x"87",x"f8",x"d0"),
  1206 => (x"05",x"a8",x"df",x"48"),
  1207 => (x"c1",x"87",x"ee",x"c1"),
  1208 => (x"c4",x"49",x"66",x"c0"),
  1209 => (x"c1",x"7e",x"69",x"81"),
  1210 => (x"6e",x"48",x"c4",x"dd"),
  1211 => (x"4a",x"a1",x"d0",x"49"),
  1212 => (x"aa",x"71",x"41",x"20"),
  1213 => (x"c1",x"87",x"f9",x"05"),
  1214 => (x"c1",x"4a",x"f1",x"c3"),
  1215 => (x"7a",x"0a",x"66",x"c0"),
  1216 => (x"66",x"c0",x"c1",x"0a"),
  1217 => (x"df",x"81",x"c9",x"49"),
  1218 => (x"66",x"c0",x"c1",x"51"),
  1219 => (x"c1",x"81",x"ca",x"49"),
  1220 => (x"c0",x"c1",x"51",x"d3"),
  1221 => (x"81",x"cb",x"49",x"66"),
  1222 => (x"c4",x"4b",x"a1",x"c4"),
  1223 => (x"78",x"6b",x"48",x"a6"),
  1224 => (x"1e",x"72",x"1e",x"71"),
  1225 => (x"48",x"d4",x"dd",x"c1"),
  1226 => (x"d0",x"49",x"66",x"cc"),
  1227 => (x"41",x"20",x"4a",x"a1"),
  1228 => (x"f9",x"05",x"aa",x"71"),
  1229 => (x"26",x"4a",x"26",x"87"),
  1230 => (x"c9",x"79",x"72",x"49"),
  1231 => (x"52",x"df",x"4a",x"a1"),
  1232 => (x"d4",x"c1",x"81",x"ca"),
  1233 => (x"48",x"a6",x"c8",x"51"),
  1234 => (x"c2",x"cf",x"78",x"c2"),
  1235 => (x"87",x"ec",x"e5",x"87"),
  1236 => (x"e5",x"87",x"ce",x"e6"),
  1237 => (x"4c",x"70",x"87",x"db"),
  1238 => (x"02",x"ac",x"fb",x"c0"),
  1239 => (x"d4",x"87",x"d0",x"c1"),
  1240 => (x"c2",x"c1",x"05",x"66"),
  1241 => (x"1e",x"1e",x"c0",x"87"),
  1242 => (x"e3",x"c1",x"1e",x"c1"),
  1243 => (x"49",x"c0",x"1e",x"c3"),
  1244 => (x"c1",x"87",x"f3",x"fb"),
  1245 => (x"c4",x"4a",x"66",x"d0"),
  1246 => (x"c7",x"49",x"6a",x"82"),
  1247 => (x"c1",x"51",x"74",x"81"),
  1248 => (x"6a",x"1e",x"d8",x"1e"),
  1249 => (x"e5",x"81",x"c8",x"49"),
  1250 => (x"86",x"d8",x"87",x"eb"),
  1251 => (x"48",x"66",x"c4",x"c1"),
  1252 => (x"c7",x"01",x"a8",x"c0"),
  1253 => (x"48",x"a6",x"c8",x"87"),
  1254 => (x"87",x"ce",x"78",x"c1"),
  1255 => (x"48",x"66",x"c4",x"c1"),
  1256 => (x"a6",x"c8",x"88",x"c1"),
  1257 => (x"e4",x"87",x"c3",x"58"),
  1258 => (x"a6",x"cc",x"87",x"f7"),
  1259 => (x"74",x"78",x"c2",x"48"),
  1260 => (x"d6",x"cd",x"02",x"9c"),
  1261 => (x"48",x"66",x"c8",x"87"),
  1262 => (x"a8",x"66",x"c8",x"c1"),
  1263 => (x"87",x"cb",x"cd",x"03"),
  1264 => (x"c0",x"48",x"a6",x"d8"),
  1265 => (x"87",x"e9",x"e3",x"78"),
  1266 => (x"d0",x"c1",x"4c",x"70"),
  1267 => (x"d6",x"c2",x"05",x"ac"),
  1268 => (x"7e",x"66",x"d8",x"87"),
  1269 => (x"70",x"87",x"cd",x"e6"),
  1270 => (x"59",x"a6",x"dc",x"49"),
  1271 => (x"70",x"87",x"d2",x"e3"),
  1272 => (x"ac",x"ec",x"c0",x"4c"),
  1273 => (x"87",x"ea",x"c1",x"05"),
  1274 => (x"cb",x"49",x"66",x"c8"),
  1275 => (x"66",x"c0",x"c1",x"91"),
  1276 => (x"4a",x"a1",x"c4",x"81"),
  1277 => (x"a1",x"c8",x"4d",x"6a"),
  1278 => (x"52",x"66",x"d8",x"4a"),
  1279 => (x"79",x"f3",x"c4",x"c1"),
  1280 => (x"70",x"87",x"ee",x"e2"),
  1281 => (x"d8",x"02",x"9c",x"4c"),
  1282 => (x"ac",x"fb",x"c0",x"87"),
  1283 => (x"74",x"87",x"d2",x"02"),
  1284 => (x"87",x"dd",x"e2",x"55"),
  1285 => (x"02",x"9c",x"4c",x"70"),
  1286 => (x"fb",x"c0",x"87",x"c7"),
  1287 => (x"ee",x"ff",x"05",x"ac"),
  1288 => (x"55",x"e0",x"c0",x"87"),
  1289 => (x"c0",x"55",x"c1",x"c2"),
  1290 => (x"66",x"d4",x"7d",x"97"),
  1291 => (x"05",x"a9",x"6e",x"49"),
  1292 => (x"66",x"c8",x"87",x"db"),
  1293 => (x"a8",x"66",x"c4",x"48"),
  1294 => (x"c8",x"87",x"ca",x"04"),
  1295 => (x"80",x"c1",x"48",x"66"),
  1296 => (x"c8",x"58",x"a6",x"cc"),
  1297 => (x"48",x"66",x"c4",x"87"),
  1298 => (x"a6",x"c8",x"88",x"c1"),
  1299 => (x"87",x"e1",x"e1",x"58"),
  1300 => (x"d0",x"c1",x"4c",x"70"),
  1301 => (x"87",x"c8",x"05",x"ac"),
  1302 => (x"c1",x"48",x"66",x"d0"),
  1303 => (x"58",x"a6",x"d4",x"80"),
  1304 => (x"02",x"ac",x"d0",x"c1"),
  1305 => (x"dc",x"87",x"ea",x"fd"),
  1306 => (x"66",x"d4",x"48",x"a6"),
  1307 => (x"48",x"66",x"d8",x"78"),
  1308 => (x"05",x"a8",x"66",x"dc"),
  1309 => (x"c0",x"87",x"e6",x"c9"),
  1310 => (x"c0",x"48",x"a6",x"e0"),
  1311 => (x"80",x"c4",x"78",x"f0"),
  1312 => (x"c4",x"78",x"66",x"cc"),
  1313 => (x"7e",x"78",x"c0",x"80"),
  1314 => (x"fb",x"c0",x"48",x"74"),
  1315 => (x"a6",x"f0",x"c0",x"88"),
  1316 => (x"02",x"98",x"70",x"58"),
  1317 => (x"48",x"87",x"e1",x"c8"),
  1318 => (x"f0",x"c0",x"88",x"cb"),
  1319 => (x"98",x"70",x"58",x"a6"),
  1320 => (x"87",x"e9",x"c0",x"02"),
  1321 => (x"c0",x"88",x"c9",x"48"),
  1322 => (x"70",x"58",x"a6",x"f0"),
  1323 => (x"e9",x"c3",x"02",x"98"),
  1324 => (x"88",x"c4",x"48",x"87"),
  1325 => (x"58",x"a6",x"f0",x"c0"),
  1326 => (x"d6",x"02",x"98",x"70"),
  1327 => (x"88",x"c1",x"48",x"87"),
  1328 => (x"58",x"a6",x"f0",x"c0"),
  1329 => (x"c3",x"02",x"98",x"70"),
  1330 => (x"e5",x"c7",x"87",x"d0"),
  1331 => (x"a6",x"e0",x"c0",x"87"),
  1332 => (x"cc",x"78",x"c0",x"48"),
  1333 => (x"80",x"c1",x"48",x"66"),
  1334 => (x"ff",x"58",x"a6",x"d0"),
  1335 => (x"70",x"87",x"d2",x"df"),
  1336 => (x"ac",x"ec",x"c0",x"4c"),
  1337 => (x"c0",x"87",x"d7",x"02"),
  1338 => (x"c0",x"02",x"66",x"e0"),
  1339 => (x"e4",x"c0",x"87",x"c7"),
  1340 => (x"c9",x"c0",x"5c",x"a6"),
  1341 => (x"c0",x"48",x"74",x"87"),
  1342 => (x"e8",x"c0",x"88",x"f0"),
  1343 => (x"ec",x"c0",x"58",x"a6"),
  1344 => (x"cd",x"c0",x"02",x"ac"),
  1345 => (x"e8",x"de",x"ff",x"87"),
  1346 => (x"c0",x"4c",x"70",x"87"),
  1347 => (x"ff",x"05",x"ac",x"ec"),
  1348 => (x"e0",x"c0",x"87",x"f3"),
  1349 => (x"66",x"d4",x"1e",x"66"),
  1350 => (x"ec",x"c0",x"1e",x"49"),
  1351 => (x"e3",x"c1",x"1e",x"66"),
  1352 => (x"66",x"d8",x"1e",x"c3"),
  1353 => (x"87",x"fe",x"f4",x"49"),
  1354 => (x"1e",x"ca",x"1e",x"c0"),
  1355 => (x"49",x"66",x"e0",x"c0"),
  1356 => (x"d8",x"c1",x"91",x"cb"),
  1357 => (x"a6",x"d8",x"81",x"66"),
  1358 => (x"78",x"a1",x"c4",x"48"),
  1359 => (x"49",x"bf",x"66",x"d8"),
  1360 => (x"87",x"f1",x"de",x"ff"),
  1361 => (x"b7",x"c0",x"86",x"d8"),
  1362 => (x"c8",x"c1",x"06",x"a8"),
  1363 => (x"de",x"1e",x"c1",x"87"),
  1364 => (x"bf",x"66",x"c8",x"1e"),
  1365 => (x"dc",x"de",x"ff",x"49"),
  1366 => (x"70",x"86",x"c8",x"87"),
  1367 => (x"08",x"c0",x"48",x"49"),
  1368 => (x"a6",x"e4",x"c0",x"88"),
  1369 => (x"a8",x"b7",x"c0",x"58"),
  1370 => (x"87",x"e9",x"c0",x"06"),
  1371 => (x"48",x"66",x"e0",x"c0"),
  1372 => (x"03",x"a8",x"b7",x"dd"),
  1373 => (x"bf",x"6e",x"87",x"df"),
  1374 => (x"66",x"e0",x"c0",x"49"),
  1375 => (x"51",x"e0",x"c0",x"81"),
  1376 => (x"81",x"c1",x"49",x"66"),
  1377 => (x"c2",x"81",x"bf",x"6e"),
  1378 => (x"e0",x"c0",x"51",x"c1"),
  1379 => (x"81",x"c2",x"49",x"66"),
  1380 => (x"c0",x"81",x"bf",x"6e"),
  1381 => (x"c4",x"7e",x"c1",x"51"),
  1382 => (x"df",x"ff",x"87",x"de"),
  1383 => (x"e4",x"c0",x"87",x"c6"),
  1384 => (x"de",x"ff",x"58",x"a6"),
  1385 => (x"e8",x"c0",x"87",x"fe"),
  1386 => (x"ec",x"c0",x"58",x"a6"),
  1387 => (x"cb",x"c0",x"05",x"a8"),
  1388 => (x"a6",x"e4",x"c0",x"87"),
  1389 => (x"66",x"e0",x"c0",x"48"),
  1390 => (x"87",x"c4",x"c0",x"78"),
  1391 => (x"87",x"f1",x"db",x"ff"),
  1392 => (x"cb",x"49",x"66",x"c8"),
  1393 => (x"66",x"c0",x"c1",x"91"),
  1394 => (x"70",x"80",x"71",x"48"),
  1395 => (x"c8",x"4a",x"6e",x"7e"),
  1396 => (x"ca",x"49",x"6e",x"82"),
  1397 => (x"66",x"e0",x"c0",x"81"),
  1398 => (x"66",x"e4",x"c0",x"51"),
  1399 => (x"c0",x"81",x"c1",x"49"),
  1400 => (x"c1",x"89",x"66",x"e0"),
  1401 => (x"70",x"30",x"71",x"48"),
  1402 => (x"71",x"89",x"c1",x"49"),
  1403 => (x"f3",x"c2",x"7a",x"97"),
  1404 => (x"c0",x"49",x"bf",x"dd"),
  1405 => (x"97",x"29",x"66",x"e0"),
  1406 => (x"71",x"48",x"4a",x"6a"),
  1407 => (x"a6",x"f0",x"c0",x"98"),
  1408 => (x"c4",x"49",x"6e",x"58"),
  1409 => (x"dc",x"4d",x"69",x"81"),
  1410 => (x"66",x"d8",x"48",x"66"),
  1411 => (x"c8",x"c0",x"02",x"a8"),
  1412 => (x"48",x"a6",x"d8",x"87"),
  1413 => (x"c5",x"c0",x"78",x"c0"),
  1414 => (x"48",x"a6",x"d8",x"87"),
  1415 => (x"66",x"d8",x"78",x"c1"),
  1416 => (x"1e",x"e0",x"c0",x"1e"),
  1417 => (x"db",x"ff",x"49",x"75"),
  1418 => (x"86",x"c8",x"87",x"cb"),
  1419 => (x"b7",x"c0",x"4c",x"70"),
  1420 => (x"d4",x"c1",x"06",x"ac"),
  1421 => (x"c0",x"85",x"74",x"87"),
  1422 => (x"89",x"74",x"49",x"e0"),
  1423 => (x"dd",x"c1",x"4b",x"75"),
  1424 => (x"fe",x"71",x"4a",x"e4"),
  1425 => (x"c2",x"87",x"fb",x"e9"),
  1426 => (x"66",x"e8",x"c0",x"85"),
  1427 => (x"c0",x"80",x"c1",x"48"),
  1428 => (x"c0",x"58",x"a6",x"ec"),
  1429 => (x"c1",x"49",x"66",x"ec"),
  1430 => (x"02",x"a9",x"70",x"81"),
  1431 => (x"d8",x"87",x"c8",x"c0"),
  1432 => (x"78",x"c0",x"48",x"a6"),
  1433 => (x"d8",x"87",x"c5",x"c0"),
  1434 => (x"78",x"c1",x"48",x"a6"),
  1435 => (x"c2",x"1e",x"66",x"d8"),
  1436 => (x"e0",x"c0",x"49",x"a4"),
  1437 => (x"70",x"88",x"71",x"48"),
  1438 => (x"49",x"75",x"1e",x"49"),
  1439 => (x"87",x"f5",x"d9",x"ff"),
  1440 => (x"b7",x"c0",x"86",x"c8"),
  1441 => (x"c0",x"ff",x"01",x"a8"),
  1442 => (x"66",x"e8",x"c0",x"87"),
  1443 => (x"87",x"d1",x"c0",x"02"),
  1444 => (x"81",x"c9",x"49",x"6e"),
  1445 => (x"51",x"66",x"e8",x"c0"),
  1446 => (x"c6",x"c1",x"48",x"6e"),
  1447 => (x"cc",x"c0",x"78",x"c3"),
  1448 => (x"c9",x"49",x"6e",x"87"),
  1449 => (x"6e",x"51",x"c2",x"81"),
  1450 => (x"f7",x"c6",x"c1",x"48"),
  1451 => (x"c0",x"7e",x"c1",x"78"),
  1452 => (x"d8",x"ff",x"87",x"c6"),
  1453 => (x"4c",x"70",x"87",x"eb"),
  1454 => (x"f5",x"c0",x"02",x"6e"),
  1455 => (x"48",x"66",x"c8",x"87"),
  1456 => (x"04",x"a8",x"66",x"c4"),
  1457 => (x"c8",x"87",x"cb",x"c0"),
  1458 => (x"80",x"c1",x"48",x"66"),
  1459 => (x"c0",x"58",x"a6",x"cc"),
  1460 => (x"66",x"c4",x"87",x"e0"),
  1461 => (x"c8",x"88",x"c1",x"48"),
  1462 => (x"d5",x"c0",x"58",x"a6"),
  1463 => (x"ac",x"c6",x"c1",x"87"),
  1464 => (x"87",x"c8",x"c0",x"05"),
  1465 => (x"c1",x"48",x"66",x"cc"),
  1466 => (x"58",x"a6",x"d0",x"80"),
  1467 => (x"87",x"f1",x"d7",x"ff"),
  1468 => (x"66",x"d0",x"4c",x"70"),
  1469 => (x"d4",x"80",x"c1",x"48"),
  1470 => (x"9c",x"74",x"58",x"a6"),
  1471 => (x"87",x"cb",x"c0",x"02"),
  1472 => (x"c1",x"48",x"66",x"c8"),
  1473 => (x"04",x"a8",x"66",x"c8"),
  1474 => (x"ff",x"87",x"f5",x"f2"),
  1475 => (x"c8",x"87",x"c9",x"d7"),
  1476 => (x"a8",x"c7",x"48",x"66"),
  1477 => (x"87",x"e5",x"c0",x"03"),
  1478 => (x"48",x"f0",x"ef",x"c2"),
  1479 => (x"66",x"c8",x"78",x"c0"),
  1480 => (x"c1",x"91",x"cb",x"49"),
  1481 => (x"c4",x"81",x"66",x"c0"),
  1482 => (x"4a",x"6a",x"4a",x"a1"),
  1483 => (x"c8",x"79",x"52",x"c0"),
  1484 => (x"80",x"c1",x"48",x"66"),
  1485 => (x"c7",x"58",x"a6",x"cc"),
  1486 => (x"db",x"ff",x"04",x"a8"),
  1487 => (x"8e",x"d0",x"ff",x"87"),
  1488 => (x"87",x"e9",x"de",x"ff"),
  1489 => (x"64",x"61",x"6f",x"4c"),
  1490 => (x"74",x"65",x"53",x"20"),
  1491 => (x"67",x"6e",x"69",x"74"),
  1492 => (x"00",x"81",x"20",x"73"),
  1493 => (x"65",x"76",x"61",x"53"),
  1494 => (x"74",x"65",x"53",x"20"),
  1495 => (x"67",x"6e",x"69",x"74"),
  1496 => (x"00",x"81",x"20",x"73"),
  1497 => (x"1e",x"00",x"20",x"3a"),
  1498 => (x"4b",x"71",x"1e",x"73"),
  1499 => (x"87",x"c6",x"02",x"9b"),
  1500 => (x"48",x"ec",x"ef",x"c2"),
  1501 => (x"1e",x"c7",x"78",x"c0"),
  1502 => (x"bf",x"ec",x"ef",x"c2"),
  1503 => (x"e1",x"c1",x"1e",x"49"),
  1504 => (x"ef",x"c2",x"1e",x"e0"),
  1505 => (x"ec",x"49",x"bf",x"e8"),
  1506 => (x"86",x"cc",x"87",x"d1"),
  1507 => (x"bf",x"e8",x"ef",x"c2"),
  1508 => (x"87",x"c7",x"e7",x"49"),
  1509 => (x"c8",x"02",x"9b",x"73"),
  1510 => (x"e0",x"e1",x"c1",x"87"),
  1511 => (x"e8",x"e5",x"c0",x"49"),
  1512 => (x"cc",x"dd",x"ff",x"87"),
  1513 => (x"f9",x"c7",x"1e",x"87"),
  1514 => (x"fe",x"49",x"c1",x"87"),
  1515 => (x"ec",x"fe",x"87",x"f9"),
  1516 => (x"98",x"70",x"87",x"d9"),
  1517 => (x"fe",x"87",x"cd",x"02"),
  1518 => (x"70",x"87",x"d6",x"f5"),
  1519 => (x"87",x"c4",x"02",x"98"),
  1520 => (x"87",x"c2",x"4a",x"c1"),
  1521 => (x"9a",x"72",x"4a",x"c0"),
  1522 => (x"c0",x"87",x"ce",x"05"),
  1523 => (x"f6",x"df",x"c1",x"1e"),
  1524 => (x"c3",x"f1",x"c0",x"49"),
  1525 => (x"fe",x"86",x"c4",x"87"),
  1526 => (x"c1",x"1e",x"c0",x"87"),
  1527 => (x"c0",x"49",x"c1",x"e0"),
  1528 => (x"c0",x"87",x"f5",x"f0"),
  1529 => (x"ca",x"c2",x"c1",x"1e"),
  1530 => (x"c0",x"49",x"70",x"87"),
  1531 => (x"c3",x"87",x"e9",x"f0"),
  1532 => (x"8e",x"f8",x"87",x"ef"),
  1533 => (x"44",x"53",x"4f",x"26"),
  1534 => (x"69",x"61",x"66",x"20"),
  1535 => (x"2e",x"64",x"65",x"6c"),
  1536 => (x"6f",x"6f",x"42",x"00"),
  1537 => (x"67",x"6e",x"69",x"74"),
  1538 => (x"00",x"2e",x"2e",x"2e"),
  1539 => (x"d4",x"e8",x"c0",x"1e"),
  1540 => (x"f6",x"f3",x"c0",x"87"),
  1541 => (x"26",x"87",x"f6",x"87"),
  1542 => (x"ef",x"c2",x"1e",x"4f"),
  1543 => (x"78",x"c0",x"48",x"ec"),
  1544 => (x"48",x"e8",x"ef",x"c2"),
  1545 => (x"fc",x"fd",x"78",x"c0"),
  1546 => (x"c0",x"87",x"e1",x"87"),
  1547 => (x"20",x"4f",x"26",x"48"),
  1548 => (x"20",x"20",x"20",x"20"),
  1549 => (x"20",x"20",x"20",x"20"),
  1550 => (x"20",x"20",x"20",x"20"),
  1551 => (x"74",x"69",x"78",x"45"),
  1552 => (x"20",x"20",x"20",x"20"),
  1553 => (x"20",x"20",x"20",x"20"),
  1554 => (x"20",x"20",x"20",x"20"),
  1555 => (x"20",x"80",x"00",x"81"),
  1556 => (x"20",x"20",x"20",x"20"),
  1557 => (x"20",x"20",x"20",x"20"),
  1558 => (x"42",x"20",x"20",x"20"),
  1559 => (x"00",x"6b",x"63",x"61"),
  1560 => (x"00",x"00",x"11",x"33"),
  1561 => (x"00",x"00",x"2c",x"01"),
  1562 => (x"33",x"00",x"00",x"00"),
  1563 => (x"1f",x"00",x"00",x"11"),
  1564 => (x"00",x"00",x"00",x"2c"),
  1565 => (x"11",x"33",x"00",x"00"),
  1566 => (x"2c",x"3d",x"00",x"00"),
  1567 => (x"00",x"00",x"00",x"00"),
  1568 => (x"00",x"11",x"33",x"00"),
  1569 => (x"00",x"2c",x"5b",x"00"),
  1570 => (x"00",x"00",x"00",x"00"),
  1571 => (x"00",x"00",x"11",x"33"),
  1572 => (x"00",x"00",x"2c",x"79"),
  1573 => (x"33",x"00",x"00",x"00"),
  1574 => (x"97",x"00",x"00",x"11"),
  1575 => (x"00",x"00",x"00",x"2c"),
  1576 => (x"11",x"33",x"00",x"00"),
  1577 => (x"2c",x"b5",x"00",x"00"),
  1578 => (x"00",x"00",x"00",x"00"),
  1579 => (x"00",x"11",x"33",x"00"),
  1580 => (x"00",x"00",x"00",x"00"),
  1581 => (x"00",x"00",x"00",x"00"),
  1582 => (x"00",x"00",x"11",x"c8"),
  1583 => (x"00",x"00",x"00",x"00"),
  1584 => (x"4c",x"00",x"00",x"00"),
  1585 => (x"20",x"64",x"61",x"6f"),
  1586 => (x"1e",x"00",x"2e",x"2a"),
  1587 => (x"c0",x"48",x"f0",x"fe"),
  1588 => (x"79",x"09",x"cd",x"78"),
  1589 => (x"1e",x"4f",x"26",x"09"),
  1590 => (x"bf",x"f0",x"fe",x"1e"),
  1591 => (x"26",x"26",x"48",x"7e"),
  1592 => (x"f0",x"fe",x"1e",x"4f"),
  1593 => (x"26",x"78",x"c1",x"48"),
  1594 => (x"f0",x"fe",x"1e",x"4f"),
  1595 => (x"26",x"78",x"c0",x"48"),
  1596 => (x"4a",x"71",x"1e",x"4f"),
  1597 => (x"26",x"52",x"52",x"c0"),
  1598 => (x"5b",x"5e",x"0e",x"4f"),
  1599 => (x"f4",x"0e",x"5d",x"5c"),
  1600 => (x"97",x"4d",x"71",x"86"),
  1601 => (x"a5",x"c1",x"7e",x"6d"),
  1602 => (x"48",x"6c",x"97",x"4c"),
  1603 => (x"6e",x"58",x"a6",x"c8"),
  1604 => (x"a8",x"66",x"c4",x"48"),
  1605 => (x"ff",x"87",x"c5",x"05"),
  1606 => (x"87",x"e6",x"c0",x"48"),
  1607 => (x"c2",x"87",x"ca",x"ff"),
  1608 => (x"6c",x"97",x"49",x"a5"),
  1609 => (x"4b",x"a3",x"71",x"4b"),
  1610 => (x"97",x"4b",x"6b",x"97"),
  1611 => (x"48",x"6e",x"7e",x"6c"),
  1612 => (x"a6",x"c8",x"80",x"c1"),
  1613 => (x"cc",x"98",x"c7",x"58"),
  1614 => (x"97",x"70",x"58",x"a6"),
  1615 => (x"87",x"e1",x"fe",x"7c"),
  1616 => (x"8e",x"f4",x"48",x"73"),
  1617 => (x"4c",x"26",x"4d",x"26"),
  1618 => (x"4f",x"26",x"4b",x"26"),
  1619 => (x"5c",x"5b",x"5e",x"0e"),
  1620 => (x"71",x"86",x"f4",x"0e"),
  1621 => (x"4a",x"66",x"d8",x"4c"),
  1622 => (x"c2",x"9a",x"ff",x"c3"),
  1623 => (x"6c",x"97",x"4b",x"a4"),
  1624 => (x"49",x"a1",x"73",x"49"),
  1625 => (x"6c",x"97",x"51",x"72"),
  1626 => (x"c1",x"48",x"6e",x"7e"),
  1627 => (x"58",x"a6",x"c8",x"80"),
  1628 => (x"a6",x"cc",x"98",x"c7"),
  1629 => (x"f4",x"54",x"70",x"58"),
  1630 => (x"87",x"ca",x"ff",x"8e"),
  1631 => (x"e8",x"fd",x"1e",x"1e"),
  1632 => (x"4a",x"bf",x"e0",x"87"),
  1633 => (x"c0",x"e0",x"c0",x"49"),
  1634 => (x"87",x"cb",x"02",x"99"),
  1635 => (x"f3",x"c2",x"1e",x"72"),
  1636 => (x"f7",x"fe",x"49",x"d3"),
  1637 => (x"fc",x"86",x"c4",x"87"),
  1638 => (x"7e",x"70",x"87",x"fd"),
  1639 => (x"26",x"87",x"c2",x"fd"),
  1640 => (x"c2",x"1e",x"4f",x"26"),
  1641 => (x"fd",x"49",x"d3",x"f3"),
  1642 => (x"e5",x"c1",x"87",x"c7"),
  1643 => (x"da",x"fc",x"49",x"fc"),
  1644 => (x"87",x"d9",x"c5",x"87"),
  1645 => (x"5e",x"0e",x"4f",x"26"),
  1646 => (x"0e",x"5d",x"5c",x"5b"),
  1647 => (x"bf",x"f2",x"f3",x"c2"),
  1648 => (x"ca",x"e8",x"c1",x"4a"),
  1649 => (x"72",x"4c",x"49",x"bf"),
  1650 => (x"fc",x"4d",x"71",x"bc"),
  1651 => (x"4b",x"c0",x"87",x"db"),
  1652 => (x"99",x"d0",x"49",x"74"),
  1653 => (x"75",x"87",x"d5",x"02"),
  1654 => (x"71",x"99",x"d0",x"49"),
  1655 => (x"c1",x"1e",x"c0",x"1e"),
  1656 => (x"73",x"4a",x"dc",x"ee"),
  1657 => (x"c0",x"49",x"12",x"82"),
  1658 => (x"86",x"c8",x"87",x"e4"),
  1659 => (x"83",x"2d",x"2c",x"c1"),
  1660 => (x"ff",x"04",x"ab",x"c8"),
  1661 => (x"e8",x"fb",x"87",x"da"),
  1662 => (x"ca",x"e8",x"c1",x"87"),
  1663 => (x"f2",x"f3",x"c2",x"48"),
  1664 => (x"4d",x"26",x"78",x"bf"),
  1665 => (x"4b",x"26",x"4c",x"26"),
  1666 => (x"00",x"00",x"4f",x"26"),
  1667 => (x"ff",x"1e",x"00",x"00"),
  1668 => (x"e1",x"c8",x"48",x"d0"),
  1669 => (x"48",x"d4",x"ff",x"78"),
  1670 => (x"66",x"c4",x"78",x"c5"),
  1671 => (x"c3",x"87",x"c3",x"02"),
  1672 => (x"66",x"c8",x"78",x"e0"),
  1673 => (x"ff",x"87",x"c6",x"02"),
  1674 => (x"f0",x"c3",x"48",x"d4"),
  1675 => (x"48",x"d4",x"ff",x"78"),
  1676 => (x"d0",x"ff",x"78",x"71"),
  1677 => (x"78",x"e1",x"c8",x"48"),
  1678 => (x"26",x"78",x"e0",x"c0"),
  1679 => (x"5b",x"5e",x"0e",x"4f"),
  1680 => (x"4c",x"71",x"0e",x"5c"),
  1681 => (x"49",x"d3",x"f3",x"c2"),
  1682 => (x"70",x"87",x"ee",x"fa"),
  1683 => (x"aa",x"b7",x"c0",x"4a"),
  1684 => (x"87",x"e3",x"c2",x"04"),
  1685 => (x"05",x"aa",x"e0",x"c3"),
  1686 => (x"ec",x"c1",x"87",x"c9"),
  1687 => (x"78",x"c1",x"48",x"c0"),
  1688 => (x"c3",x"87",x"d4",x"c2"),
  1689 => (x"c9",x"05",x"aa",x"f0"),
  1690 => (x"fc",x"eb",x"c1",x"87"),
  1691 => (x"c1",x"78",x"c1",x"48"),
  1692 => (x"ec",x"c1",x"87",x"f5"),
  1693 => (x"c7",x"02",x"bf",x"c0"),
  1694 => (x"c2",x"4b",x"72",x"87"),
  1695 => (x"87",x"c2",x"b3",x"c0"),
  1696 => (x"9c",x"74",x"4b",x"72"),
  1697 => (x"c1",x"87",x"d1",x"05"),
  1698 => (x"1e",x"bf",x"fc",x"eb"),
  1699 => (x"bf",x"c0",x"ec",x"c1"),
  1700 => (x"fd",x"49",x"72",x"1e"),
  1701 => (x"86",x"c8",x"87",x"f8"),
  1702 => (x"bf",x"fc",x"eb",x"c1"),
  1703 => (x"87",x"e0",x"c0",x"02"),
  1704 => (x"b7",x"c4",x"49",x"73"),
  1705 => (x"ed",x"c1",x"91",x"29"),
  1706 => (x"4a",x"73",x"81",x"dc"),
  1707 => (x"92",x"c2",x"9a",x"cf"),
  1708 => (x"30",x"72",x"48",x"c1"),
  1709 => (x"ba",x"ff",x"4a",x"70"),
  1710 => (x"98",x"69",x"48",x"72"),
  1711 => (x"87",x"db",x"79",x"70"),
  1712 => (x"b7",x"c4",x"49",x"73"),
  1713 => (x"ed",x"c1",x"91",x"29"),
  1714 => (x"4a",x"73",x"81",x"dc"),
  1715 => (x"92",x"c2",x"9a",x"cf"),
  1716 => (x"30",x"72",x"48",x"c3"),
  1717 => (x"69",x"48",x"4a",x"70"),
  1718 => (x"c1",x"79",x"70",x"b0"),
  1719 => (x"c0",x"48",x"c0",x"ec"),
  1720 => (x"fc",x"eb",x"c1",x"78"),
  1721 => (x"c2",x"78",x"c0",x"48"),
  1722 => (x"f8",x"49",x"d3",x"f3"),
  1723 => (x"4a",x"70",x"87",x"cb"),
  1724 => (x"03",x"aa",x"b7",x"c0"),
  1725 => (x"c0",x"87",x"dd",x"fd"),
  1726 => (x"87",x"c8",x"fc",x"48"),
  1727 => (x"00",x"00",x"00",x"00"),
  1728 => (x"00",x"00",x"00",x"00"),
  1729 => (x"49",x"4a",x"71",x"1e"),
  1730 => (x"26",x"87",x"f2",x"fc"),
  1731 => (x"4a",x"c0",x"1e",x"4f"),
  1732 => (x"91",x"c4",x"49",x"72"),
  1733 => (x"81",x"dc",x"ed",x"c1"),
  1734 => (x"82",x"c1",x"79",x"c0"),
  1735 => (x"04",x"aa",x"b7",x"d0"),
  1736 => (x"4f",x"26",x"87",x"ee"),
  1737 => (x"5c",x"5b",x"5e",x"0e"),
  1738 => (x"4d",x"71",x"0e",x"5d"),
  1739 => (x"75",x"87",x"fa",x"f6"),
  1740 => (x"2a",x"b7",x"c4",x"4a"),
  1741 => (x"dc",x"ed",x"c1",x"92"),
  1742 => (x"cf",x"4c",x"75",x"82"),
  1743 => (x"6a",x"94",x"c2",x"9c"),
  1744 => (x"2b",x"74",x"4b",x"49"),
  1745 => (x"48",x"c2",x"9b",x"c3"),
  1746 => (x"4c",x"70",x"30",x"74"),
  1747 => (x"48",x"74",x"bc",x"ff"),
  1748 => (x"7a",x"70",x"98",x"71"),
  1749 => (x"73",x"87",x"ca",x"f6"),
  1750 => (x"87",x"e6",x"fa",x"48"),
  1751 => (x"00",x"00",x"00",x"00"),
  1752 => (x"00",x"00",x"00",x"00"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"00",x"00",x"00"),
  1755 => (x"00",x"00",x"00",x"00"),
  1756 => (x"00",x"00",x"00",x"00"),
  1757 => (x"00",x"00",x"00",x"00"),
  1758 => (x"00",x"00",x"00",x"00"),
  1759 => (x"00",x"00",x"00",x"00"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"25",x"26",x"1e",x"16"),
  1768 => (x"3e",x"3d",x"36",x"2e"),
  1769 => (x"48",x"d0",x"ff",x"1e"),
  1770 => (x"71",x"78",x"e1",x"c8"),
  1771 => (x"08",x"d4",x"ff",x"48"),
  1772 => (x"1e",x"4f",x"26",x"78"),
  1773 => (x"c8",x"48",x"d0",x"ff"),
  1774 => (x"48",x"71",x"78",x"e1"),
  1775 => (x"78",x"08",x"d4",x"ff"),
  1776 => (x"ff",x"48",x"66",x"c4"),
  1777 => (x"26",x"78",x"08",x"d4"),
  1778 => (x"4a",x"71",x"1e",x"4f"),
  1779 => (x"1e",x"49",x"66",x"c4"),
  1780 => (x"de",x"ff",x"49",x"72"),
  1781 => (x"48",x"d0",x"ff",x"87"),
  1782 => (x"26",x"78",x"e0",x"c0"),
  1783 => (x"71",x"1e",x"4f",x"26"),
  1784 => (x"aa",x"b7",x"c2",x"4a"),
  1785 => (x"82",x"87",x"c3",x"03"),
  1786 => (x"82",x"ce",x"87",x"c2"),
  1787 => (x"72",x"1e",x"66",x"c4"),
  1788 => (x"87",x"d5",x"ff",x"49"),
  1789 => (x"1e",x"4f",x"26",x"26"),
  1790 => (x"c3",x"4a",x"d4",x"ff"),
  1791 => (x"d0",x"ff",x"7a",x"ff"),
  1792 => (x"78",x"e1",x"c8",x"48"),
  1793 => (x"f3",x"c2",x"7a",x"de"),
  1794 => (x"49",x"7a",x"bf",x"dd"),
  1795 => (x"70",x"28",x"c8",x"48"),
  1796 => (x"d0",x"48",x"71",x"7a"),
  1797 => (x"71",x"7a",x"70",x"28"),
  1798 => (x"70",x"28",x"d8",x"48"),
  1799 => (x"48",x"d0",x"ff",x"7a"),
  1800 => (x"26",x"78",x"e0",x"c0"),
  1801 => (x"5b",x"5e",x"0e",x"4f"),
  1802 => (x"71",x"0e",x"5d",x"5c"),
  1803 => (x"dd",x"f3",x"c2",x"4c"),
  1804 => (x"74",x"4b",x"4d",x"bf"),
  1805 => (x"9b",x"66",x"d0",x"2b"),
  1806 => (x"66",x"d4",x"83",x"c1"),
  1807 => (x"87",x"c2",x"04",x"ab"),
  1808 => (x"4a",x"74",x"4b",x"c0"),
  1809 => (x"72",x"49",x"66",x"d0"),
  1810 => (x"75",x"b9",x"ff",x"31"),
  1811 => (x"72",x"48",x"73",x"99"),
  1812 => (x"48",x"4a",x"70",x"30"),
  1813 => (x"f3",x"c2",x"b0",x"71"),
  1814 => (x"da",x"fe",x"58",x"e1"),
  1815 => (x"26",x"4d",x"26",x"87"),
  1816 => (x"26",x"4b",x"26",x"4c"),
  1817 => (x"d0",x"ff",x"1e",x"4f"),
  1818 => (x"78",x"c9",x"c8",x"48"),
  1819 => (x"d4",x"ff",x"48",x"71"),
  1820 => (x"4f",x"26",x"78",x"08"),
  1821 => (x"49",x"4a",x"71",x"1e"),
  1822 => (x"d0",x"ff",x"87",x"eb"),
  1823 => (x"26",x"78",x"c8",x"48"),
  1824 => (x"1e",x"73",x"1e",x"4f"),
  1825 => (x"f3",x"c2",x"4b",x"71"),
  1826 => (x"c3",x"02",x"bf",x"ed"),
  1827 => (x"87",x"eb",x"c2",x"87"),
  1828 => (x"c8",x"48",x"d0",x"ff"),
  1829 => (x"49",x"73",x"78",x"c9"),
  1830 => (x"ff",x"b1",x"e0",x"c0"),
  1831 => (x"78",x"71",x"48",x"d4"),
  1832 => (x"48",x"e1",x"f3",x"c2"),
  1833 => (x"66",x"c8",x"78",x"c0"),
  1834 => (x"c3",x"87",x"c5",x"02"),
  1835 => (x"87",x"c2",x"49",x"ff"),
  1836 => (x"f3",x"c2",x"49",x"c0"),
  1837 => (x"66",x"cc",x"59",x"e9"),
  1838 => (x"c5",x"87",x"c6",x"02"),
  1839 => (x"c4",x"4a",x"d5",x"d5"),
  1840 => (x"ff",x"ff",x"cf",x"87"),
  1841 => (x"ed",x"f3",x"c2",x"4a"),
  1842 => (x"ed",x"f3",x"c2",x"5a"),
  1843 => (x"c4",x"78",x"c1",x"48"),
  1844 => (x"26",x"4d",x"26",x"87"),
  1845 => (x"26",x"4b",x"26",x"4c"),
  1846 => (x"5b",x"5e",x"0e",x"4f"),
  1847 => (x"71",x"0e",x"5d",x"5c"),
  1848 => (x"e9",x"f3",x"c2",x"4a"),
  1849 => (x"9a",x"72",x"4c",x"bf"),
  1850 => (x"49",x"87",x"cb",x"02"),
  1851 => (x"f1",x"c1",x"91",x"c8"),
  1852 => (x"83",x"71",x"4b",x"f7"),
  1853 => (x"f5",x"c1",x"87",x"c4"),
  1854 => (x"4d",x"c0",x"4b",x"f7"),
  1855 => (x"99",x"74",x"49",x"13"),
  1856 => (x"bf",x"e5",x"f3",x"c2"),
  1857 => (x"48",x"d4",x"ff",x"b9"),
  1858 => (x"b7",x"c1",x"78",x"71"),
  1859 => (x"b7",x"c8",x"85",x"2c"),
  1860 => (x"87",x"e8",x"04",x"ad"),
  1861 => (x"bf",x"e1",x"f3",x"c2"),
  1862 => (x"c2",x"80",x"c8",x"48"),
  1863 => (x"fe",x"58",x"e5",x"f3"),
  1864 => (x"73",x"1e",x"87",x"ef"),
  1865 => (x"13",x"4b",x"71",x"1e"),
  1866 => (x"cb",x"02",x"9a",x"4a"),
  1867 => (x"fe",x"49",x"72",x"87"),
  1868 => (x"4a",x"13",x"87",x"e7"),
  1869 => (x"87",x"f5",x"05",x"9a"),
  1870 => (x"1e",x"87",x"da",x"fe"),
  1871 => (x"bf",x"e1",x"f3",x"c2"),
  1872 => (x"e1",x"f3",x"c2",x"49"),
  1873 => (x"78",x"a1",x"c1",x"48"),
  1874 => (x"a9",x"b7",x"c0",x"c4"),
  1875 => (x"ff",x"87",x"db",x"03"),
  1876 => (x"f3",x"c2",x"48",x"d4"),
  1877 => (x"c2",x"78",x"bf",x"e5"),
  1878 => (x"49",x"bf",x"e1",x"f3"),
  1879 => (x"48",x"e1",x"f3",x"c2"),
  1880 => (x"c4",x"78",x"a1",x"c1"),
  1881 => (x"04",x"a9",x"b7",x"c0"),
  1882 => (x"d0",x"ff",x"87",x"e5"),
  1883 => (x"c2",x"78",x"c8",x"48"),
  1884 => (x"c0",x"48",x"ed",x"f3"),
  1885 => (x"00",x"4f",x"26",x"78"),
  1886 => (x"00",x"00",x"00",x"00"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"5f",x"5f",x"00",x"00"),
  1889 => (x"00",x"00",x"00",x"00"),
  1890 => (x"03",x"00",x"03",x"03"),
  1891 => (x"14",x"00",x"00",x"03"),
  1892 => (x"7f",x"14",x"7f",x"7f"),
  1893 => (x"00",x"00",x"14",x"7f"),
  1894 => (x"6b",x"6b",x"2e",x"24"),
  1895 => (x"4c",x"00",x"12",x"3a"),
  1896 => (x"6c",x"18",x"36",x"6a"),
  1897 => (x"30",x"00",x"32",x"56"),
  1898 => (x"77",x"59",x"4f",x"7e"),
  1899 => (x"00",x"40",x"68",x"3a"),
  1900 => (x"03",x"07",x"04",x"00"),
  1901 => (x"00",x"00",x"00",x"00"),
  1902 => (x"63",x"3e",x"1c",x"00"),
  1903 => (x"00",x"00",x"00",x"41"),
  1904 => (x"3e",x"63",x"41",x"00"),
  1905 => (x"08",x"00",x"00",x"1c"),
  1906 => (x"1c",x"1c",x"3e",x"2a"),
  1907 => (x"00",x"08",x"2a",x"3e"),
  1908 => (x"3e",x"3e",x"08",x"08"),
  1909 => (x"00",x"00",x"08",x"08"),
  1910 => (x"60",x"e0",x"80",x"00"),
  1911 => (x"00",x"00",x"00",x"00"),
  1912 => (x"08",x"08",x"08",x"08"),
  1913 => (x"00",x"00",x"08",x"08"),
  1914 => (x"60",x"60",x"00",x"00"),
  1915 => (x"40",x"00",x"00",x"00"),
  1916 => (x"0c",x"18",x"30",x"60"),
  1917 => (x"00",x"01",x"03",x"06"),
  1918 => (x"4d",x"59",x"7f",x"3e"),
  1919 => (x"00",x"00",x"3e",x"7f"),
  1920 => (x"7f",x"7f",x"06",x"04"),
  1921 => (x"00",x"00",x"00",x"00"),
  1922 => (x"59",x"71",x"63",x"42"),
  1923 => (x"00",x"00",x"46",x"4f"),
  1924 => (x"49",x"49",x"63",x"22"),
  1925 => (x"18",x"00",x"36",x"7f"),
  1926 => (x"7f",x"13",x"16",x"1c"),
  1927 => (x"00",x"00",x"10",x"7f"),
  1928 => (x"45",x"45",x"67",x"27"),
  1929 => (x"00",x"00",x"39",x"7d"),
  1930 => (x"49",x"4b",x"7e",x"3c"),
  1931 => (x"00",x"00",x"30",x"79"),
  1932 => (x"79",x"71",x"01",x"01"),
  1933 => (x"00",x"00",x"07",x"0f"),
  1934 => (x"49",x"49",x"7f",x"36"),
  1935 => (x"00",x"00",x"36",x"7f"),
  1936 => (x"69",x"49",x"4f",x"06"),
  1937 => (x"00",x"00",x"1e",x"3f"),
  1938 => (x"66",x"66",x"00",x"00"),
  1939 => (x"00",x"00",x"00",x"00"),
  1940 => (x"66",x"e6",x"80",x"00"),
  1941 => (x"00",x"00",x"00",x"00"),
  1942 => (x"14",x"14",x"08",x"08"),
  1943 => (x"00",x"00",x"22",x"22"),
  1944 => (x"14",x"14",x"14",x"14"),
  1945 => (x"00",x"00",x"14",x"14"),
  1946 => (x"14",x"14",x"22",x"22"),
  1947 => (x"00",x"00",x"08",x"08"),
  1948 => (x"59",x"51",x"03",x"02"),
  1949 => (x"3e",x"00",x"06",x"0f"),
  1950 => (x"55",x"5d",x"41",x"7f"),
  1951 => (x"00",x"00",x"1e",x"1f"),
  1952 => (x"09",x"09",x"7f",x"7e"),
  1953 => (x"00",x"00",x"7e",x"7f"),
  1954 => (x"49",x"49",x"7f",x"7f"),
  1955 => (x"00",x"00",x"36",x"7f"),
  1956 => (x"41",x"63",x"3e",x"1c"),
  1957 => (x"00",x"00",x"41",x"41"),
  1958 => (x"63",x"41",x"7f",x"7f"),
  1959 => (x"00",x"00",x"1c",x"3e"),
  1960 => (x"49",x"49",x"7f",x"7f"),
  1961 => (x"00",x"00",x"41",x"41"),
  1962 => (x"09",x"09",x"7f",x"7f"),
  1963 => (x"00",x"00",x"01",x"01"),
  1964 => (x"49",x"41",x"7f",x"3e"),
  1965 => (x"00",x"00",x"7a",x"7b"),
  1966 => (x"08",x"08",x"7f",x"7f"),
  1967 => (x"00",x"00",x"7f",x"7f"),
  1968 => (x"7f",x"7f",x"41",x"00"),
  1969 => (x"00",x"00",x"00",x"41"),
  1970 => (x"40",x"40",x"60",x"20"),
  1971 => (x"7f",x"00",x"3f",x"7f"),
  1972 => (x"36",x"1c",x"08",x"7f"),
  1973 => (x"00",x"00",x"41",x"63"),
  1974 => (x"40",x"40",x"7f",x"7f"),
  1975 => (x"7f",x"00",x"40",x"40"),
  1976 => (x"06",x"0c",x"06",x"7f"),
  1977 => (x"7f",x"00",x"7f",x"7f"),
  1978 => (x"18",x"0c",x"06",x"7f"),
  1979 => (x"00",x"00",x"7f",x"7f"),
  1980 => (x"41",x"41",x"7f",x"3e"),
  1981 => (x"00",x"00",x"3e",x"7f"),
  1982 => (x"09",x"09",x"7f",x"7f"),
  1983 => (x"3e",x"00",x"06",x"0f"),
  1984 => (x"7f",x"61",x"41",x"7f"),
  1985 => (x"00",x"00",x"40",x"7e"),
  1986 => (x"19",x"09",x"7f",x"7f"),
  1987 => (x"00",x"00",x"66",x"7f"),
  1988 => (x"59",x"4d",x"6f",x"26"),
  1989 => (x"00",x"00",x"32",x"7b"),
  1990 => (x"7f",x"7f",x"01",x"01"),
  1991 => (x"00",x"00",x"01",x"01"),
  1992 => (x"40",x"40",x"7f",x"3f"),
  1993 => (x"00",x"00",x"3f",x"7f"),
  1994 => (x"70",x"70",x"3f",x"0f"),
  1995 => (x"7f",x"00",x"0f",x"3f"),
  1996 => (x"30",x"18",x"30",x"7f"),
  1997 => (x"41",x"00",x"7f",x"7f"),
  1998 => (x"1c",x"1c",x"36",x"63"),
  1999 => (x"01",x"41",x"63",x"36"),
  2000 => (x"7c",x"7c",x"06",x"03"),
  2001 => (x"61",x"01",x"03",x"06"),
  2002 => (x"47",x"4d",x"59",x"71"),
  2003 => (x"00",x"00",x"41",x"43"),
  2004 => (x"41",x"7f",x"7f",x"00"),
  2005 => (x"01",x"00",x"00",x"41"),
  2006 => (x"18",x"0c",x"06",x"03"),
  2007 => (x"00",x"40",x"60",x"30"),
  2008 => (x"7f",x"41",x"41",x"00"),
  2009 => (x"08",x"00",x"00",x"7f"),
  2010 => (x"06",x"03",x"06",x"0c"),
  2011 => (x"80",x"00",x"08",x"0c"),
  2012 => (x"80",x"80",x"80",x"80"),
  2013 => (x"00",x"00",x"80",x"80"),
  2014 => (x"07",x"03",x"00",x"00"),
  2015 => (x"00",x"00",x"00",x"04"),
  2016 => (x"54",x"54",x"74",x"20"),
  2017 => (x"00",x"00",x"78",x"7c"),
  2018 => (x"44",x"44",x"7f",x"7f"),
  2019 => (x"00",x"00",x"38",x"7c"),
  2020 => (x"44",x"44",x"7c",x"38"),
  2021 => (x"00",x"00",x"00",x"44"),
  2022 => (x"44",x"44",x"7c",x"38"),
  2023 => (x"00",x"00",x"7f",x"7f"),
  2024 => (x"54",x"54",x"7c",x"38"),
  2025 => (x"00",x"00",x"18",x"5c"),
  2026 => (x"05",x"7f",x"7e",x"04"),
  2027 => (x"00",x"00",x"00",x"05"),
  2028 => (x"a4",x"a4",x"bc",x"18"),
  2029 => (x"00",x"00",x"7c",x"fc"),
  2030 => (x"04",x"04",x"7f",x"7f"),
  2031 => (x"00",x"00",x"78",x"7c"),
  2032 => (x"7d",x"3d",x"00",x"00"),
  2033 => (x"00",x"00",x"00",x"40"),
  2034 => (x"fd",x"80",x"80",x"80"),
  2035 => (x"00",x"00",x"00",x"7d"),
  2036 => (x"38",x"10",x"7f",x"7f"),
  2037 => (x"00",x"00",x"44",x"6c"),
  2038 => (x"7f",x"3f",x"00",x"00"),
  2039 => (x"7c",x"00",x"00",x"40"),
  2040 => (x"0c",x"18",x"0c",x"7c"),
  2041 => (x"00",x"00",x"78",x"7c"),
  2042 => (x"04",x"04",x"7c",x"7c"),
  2043 => (x"00",x"00",x"78",x"7c"),
  2044 => (x"44",x"44",x"7c",x"38"),
  2045 => (x"00",x"00",x"38",x"7c"),
  2046 => (x"24",x"24",x"fc",x"fc"),
  2047 => (x"00",x"00",x"18",x"3c"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

