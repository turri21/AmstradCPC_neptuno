library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"24243c18",
     1 => x"0000fcfc",
     2 => x"04047c7c",
     3 => x"0000080c",
     4 => x"54545c48",
     5 => x"00002074",
     6 => x"447f3f04",
     7 => x"00000044",
     8 => x"40407c3c",
     9 => x"00007c7c",
    10 => x"60603c1c",
    11 => x"3c001c3c",
    12 => x"6030607c",
    13 => x"44003c7c",
    14 => x"3810386c",
    15 => x"0000446c",
    16 => x"60e0bc1c",
    17 => x"00001c3c",
    18 => x"5c746444",
    19 => x"0000444c",
    20 => x"773e0808",
    21 => x"00004141",
    22 => x"7f7f0000",
    23 => x"00000000",
    24 => x"3e774141",
    25 => x"02000808",
    26 => x"02030101",
    27 => x"7f000102",
    28 => x"7f7f7f7f",
    29 => x"08007f7f",
    30 => x"3e1c1c08",
    31 => x"7f7f7f3e",
    32 => x"1c3e3e7f",
    33 => x"0008081c",
    34 => x"7c7c1810",
    35 => x"00001018",
    36 => x"7c7c3010",
    37 => x"10001030",
    38 => x"78606030",
    39 => x"4200061e",
    40 => x"3c183c66",
    41 => x"78004266",
    42 => x"c6c26a38",
    43 => x"6000386c",
    44 => x"00600000",
    45 => x"0e006000",
    46 => x"5d5c5b5e",
    47 => x"4c711e0e",
    48 => x"bffef3c2",
    49 => x"c04bc04d",
    50 => x"02ab741e",
    51 => x"a6c487c7",
    52 => x"c578c048",
    53 => x"48a6c487",
    54 => x"66c478c1",
    55 => x"ee49731e",
    56 => x"86c887df",
    57 => x"ef49e0c0",
    58 => x"a5c487ef",
    59 => x"f0496a4a",
    60 => x"c6f187f0",
    61 => x"c185cb87",
    62 => x"abb7c883",
    63 => x"87c7ff04",
    64 => x"264d2626",
    65 => x"264b264c",
    66 => x"4a711e4f",
    67 => x"5ac2f4c2",
    68 => x"48c2f4c2",
    69 => x"fe4978c7",
    70 => x"4f2687dd",
    71 => x"711e731e",
    72 => x"aab7c04a",
    73 => x"c287d303",
    74 => x"05bfedd1",
    75 => x"4bc187c4",
    76 => x"4bc087c2",
    77 => x"5bf1d1c2",
    78 => x"d1c287c4",
    79 => x"d1c25af1",
    80 => x"c14abfed",
    81 => x"a2c0c19a",
    82 => x"87e8ec49",
    83 => x"d1c248fc",
    84 => x"fe78bfed",
    85 => x"711e87ef",
    86 => x"1e66c44a",
    87 => x"fde94972",
    88 => x"4f262687",
    89 => x"edd1c21e",
    90 => x"d7e649bf",
    91 => x"f6f3c287",
    92 => x"78bfe848",
    93 => x"48f2f3c2",
    94 => x"c278bfec",
    95 => x"4abff6f3",
    96 => x"99ffc349",
    97 => x"722ab7c8",
    98 => x"c2b07148",
    99 => x"2658fef3",
   100 => x"5b5e0e4f",
   101 => x"710e5d5c",
   102 => x"87c8ff4b",
   103 => x"48f1f3c2",
   104 => x"497350c0",
   105 => x"7087fde5",
   106 => x"9cc24c49",
   107 => x"cb49eecb",
   108 => x"497087c3",
   109 => x"f1f3c24d",
   110 => x"c105bf97",
   111 => x"66d087e2",
   112 => x"faf3c249",
   113 => x"d60599bf",
   114 => x"4966d487",
   115 => x"bff2f3c2",
   116 => x"87cb0599",
   117 => x"cbe54973",
   118 => x"02987087",
   119 => x"c187c1c1",
   120 => x"87c0fe4c",
   121 => x"d8ca4975",
   122 => x"02987087",
   123 => x"f3c287c6",
   124 => x"50c148f1",
   125 => x"97f1f3c2",
   126 => x"e3c005bf",
   127 => x"faf3c287",
   128 => x"66d049bf",
   129 => x"d6ff0599",
   130 => x"f2f3c287",
   131 => x"66d449bf",
   132 => x"caff0599",
   133 => x"e4497387",
   134 => x"987087ca",
   135 => x"87fffe05",
   136 => x"dcfb4874",
   137 => x"5b5e0e87",
   138 => x"f40e5d5c",
   139 => x"4c4dc086",
   140 => x"c47ebfec",
   141 => x"f3c248a6",
   142 => x"c178bffe",
   143 => x"c71ec01e",
   144 => x"87cdfd49",
   145 => x"987086c8",
   146 => x"ff87cd02",
   147 => x"87ccfb49",
   148 => x"e349dac1",
   149 => x"4dc187ce",
   150 => x"97f1f3c2",
   151 => x"87c302bf",
   152 => x"c287cad5",
   153 => x"4bbff6f3",
   154 => x"bfedd1c2",
   155 => x"87e9c005",
   156 => x"e249fdc3",
   157 => x"fac387ee",
   158 => x"87e8e249",
   159 => x"ffc34973",
   160 => x"c01e7199",
   161 => x"87cefb49",
   162 => x"b7c84973",
   163 => x"c11e7129",
   164 => x"87c2fb49",
   165 => x"fac586c8",
   166 => x"faf3c287",
   167 => x"029b4bbf",
   168 => x"d1c287dd",
   169 => x"c749bfe9",
   170 => x"987087d7",
   171 => x"c087c405",
   172 => x"c287d24b",
   173 => x"fcc649e0",
   174 => x"edd1c287",
   175 => x"c287c658",
   176 => x"c048e9d1",
   177 => x"c2497378",
   178 => x"87cd0599",
   179 => x"e149ebc3",
   180 => x"497087d2",
   181 => x"c20299c2",
   182 => x"734cfb87",
   183 => x"0599c149",
   184 => x"f4c387cd",
   185 => x"87fce049",
   186 => x"99c24970",
   187 => x"fa87c202",
   188 => x"c849734c",
   189 => x"87cd0599",
   190 => x"e049f5c3",
   191 => x"497087e6",
   192 => x"d40299c2",
   193 => x"c2f4c287",
   194 => x"87c902bf",
   195 => x"c288c148",
   196 => x"c258c6f4",
   197 => x"c14cff87",
   198 => x"c449734d",
   199 => x"87ce0599",
   200 => x"ff49f2c3",
   201 => x"7087fddf",
   202 => x"0299c249",
   203 => x"f4c287db",
   204 => x"487ebfc2",
   205 => x"03a8b7c7",
   206 => x"486e87cb",
   207 => x"f4c280c1",
   208 => x"c2c058c6",
   209 => x"c14cfe87",
   210 => x"49fdc34d",
   211 => x"87d4dfff",
   212 => x"99c24970",
   213 => x"c287d502",
   214 => x"02bfc2f4",
   215 => x"c287c9c0",
   216 => x"c048c2f4",
   217 => x"87c2c078",
   218 => x"4dc14cfd",
   219 => x"ff49fac3",
   220 => x"7087f1de",
   221 => x"0299c249",
   222 => x"f4c287d9",
   223 => x"c748bfc2",
   224 => x"c003a8b7",
   225 => x"f4c287c9",
   226 => x"78c748c2",
   227 => x"fc87c2c0",
   228 => x"c04dc14c",
   229 => x"c003acb7",
   230 => x"66c487d1",
   231 => x"82d8c14a",
   232 => x"c6c0026a",
   233 => x"744b6a87",
   234 => x"c00f7349",
   235 => x"1ef0c31e",
   236 => x"f749dac1",
   237 => x"86c887db",
   238 => x"c0029870",
   239 => x"a6c887e2",
   240 => x"c2f4c248",
   241 => x"66c878bf",
   242 => x"c491cb49",
   243 => x"80714866",
   244 => x"bf6e7e70",
   245 => x"87c8c002",
   246 => x"c84bbf6e",
   247 => x"0f734966",
   248 => x"c0029d75",
   249 => x"f4c287c8",
   250 => x"f349bfc2",
   251 => x"d1c287c9",
   252 => x"c002bff1",
   253 => x"c24987dd",
   254 => x"987087c7",
   255 => x"87d3c002",
   256 => x"bfc2f4c2",
   257 => x"87eff249",
   258 => x"cff449c0",
   259 => x"f1d1c287",
   260 => x"f478c048",
   261 => x"87e9f38e",
   262 => x"5c5b5e0e",
   263 => x"711e0e5d",
   264 => x"fef3c24c",
   265 => x"cdc149bf",
   266 => x"d1c14da1",
   267 => x"747e6981",
   268 => x"87cf029c",
   269 => x"744ba5c4",
   270 => x"fef3c27b",
   271 => x"c8f349bf",
   272 => x"747b6e87",
   273 => x"87c4059c",
   274 => x"87c24bc0",
   275 => x"49734bc1",
   276 => x"d487c9f3",
   277 => x"87c70266",
   278 => x"7087da49",
   279 => x"c087c24a",
   280 => x"f5d1c24a",
   281 => x"d8f2265a",
   282 => x"00000087",
   283 => x"00000000",
   284 => x"00000000",
   285 => x"4a711e00",
   286 => x"49bfc8ff",
   287 => x"2648a172",
   288 => x"c8ff1e4f",
   289 => x"c0fe89bf",
   290 => x"c0c0c0c0",
   291 => x"87c401a9",
   292 => x"87c24ac0",
   293 => x"48724ac1",
   294 => x"5e0e4f26",
   295 => x"0e5d5c5b",
   296 => x"d4ff4b71",
   297 => x"4866d04c",
   298 => x"49d678c0",
   299 => x"87f4dbff",
   300 => x"6c7cffc3",
   301 => x"99ffc349",
   302 => x"c3494d71",
   303 => x"e0c199f0",
   304 => x"87cb05a9",
   305 => x"6c7cffc3",
   306 => x"d098c348",
   307 => x"c3780866",
   308 => x"4a6c7cff",
   309 => x"c331c849",
   310 => x"4a6c7cff",
   311 => x"4972b271",
   312 => x"ffc331c8",
   313 => x"714a6c7c",
   314 => x"c84972b2",
   315 => x"7cffc331",
   316 => x"b2714a6c",
   317 => x"c048d0ff",
   318 => x"9b7378e0",
   319 => x"7287c202",
   320 => x"2648757b",
   321 => x"264c264d",
   322 => x"1e4f264b",
   323 => x"86f81e73",
   324 => x"a6c81e76",
   325 => x"87c2fe49",
   326 => x"4b7086c4",
   327 => x"a8c4486e",
   328 => x"87efc203",
   329 => x"f0c34a73",
   330 => x"aad0c19a",
   331 => x"c187c702",
   332 => x"c205aae0",
   333 => x"9bc387dd",
   334 => x"c487d802",
   335 => x"31c94966",
   336 => x"66c41e71",
   337 => x"c292d44a",
   338 => x"7249c6f4",
   339 => x"eed1fe81",
   340 => x"c286c487",
   341 => x"f6c005ab",
   342 => x"1e496e87",
   343 => x"ff49e3c0",
   344 => x"d887e6d9",
   345 => x"fbd8ff49",
   346 => x"1ec0c887",
   347 => x"49f6e2c2",
   348 => x"87fcedfd",
   349 => x"c048d0ff",
   350 => x"e2c278e0",
   351 => x"66cc1ef6",
   352 => x"c292d44a",
   353 => x"7249c6f4",
   354 => x"efcffe81",
   355 => x"c186cc87",
   356 => x"fec005ab",
   357 => x"49f2c187",
   358 => x"87f3eafd",
   359 => x"1ef6e2c2",
   360 => x"d44a66c4",
   361 => x"c6f4c292",
   362 => x"fe817249",
   363 => x"c487cace",
   364 => x"c01e4966",
   365 => x"d8ff49e3",
   366 => x"49d787cf",
   367 => x"87e4d7ff",
   368 => x"c21ec0c8",
   369 => x"fd49f6e2",
   370 => x"cc87d4ec",
   371 => x"48d0ff86",
   372 => x"f878e0c0",
   373 => x"87effc8e",
   374 => x"5c5b5e0e",
   375 => x"711e0e5d",
   376 => x"4cd4ff4d",
   377 => x"487e66d4",
   378 => x"06a8b7c4",
   379 => x"48c087c5",
   380 => x"7587e6c1",
   381 => x"d7defe49",
   382 => x"c41e7587",
   383 => x"93d44b66",
   384 => x"83c6f4c2",
   385 => x"c9fe4973",
   386 => x"83c887d3",
   387 => x"d0ff4b6b",
   388 => x"78e1c848",
   389 => x"48737cdd",
   390 => x"7098ffc3",
   391 => x"c849737c",
   392 => x"c3487129",
   393 => x"7c7098ff",
   394 => x"29d04973",
   395 => x"ffc34871",
   396 => x"737c7098",
   397 => x"7028d848",
   398 => x"7c7cc07c",
   399 => x"7c7c7c7c",
   400 => x"7c7c7c7c",
   401 => x"d0ff7c7c",
   402 => x"78e0c048",
   403 => x"dc1e66c4",
   404 => x"f4d5ff49",
   405 => x"7386c887",
   406 => x"e6fa2648",
   407 => x"5b5e0e87",
   408 => x"1e0e5d5c",
   409 => x"d4ff7e71",
   410 => x"c21e6e4b",
   411 => x"fe49d6f5",
   412 => x"c487eac7",
   413 => x"9d4d7086",
   414 => x"87c3c302",
   415 => x"bfdef5c2",
   416 => x"fe496e4c",
   417 => x"ff87c9dc",
   418 => x"c5c848d0",
   419 => x"7bd6c178",
   420 => x"7b154ac0",
   421 => x"e0c082c1",
   422 => x"f504aab7",
   423 => x"48d0ff87",
   424 => x"c5c878c4",
   425 => x"7bd3c178",
   426 => x"78c47bc1",
   427 => x"c1029c74",
   428 => x"e2c287fc",
   429 => x"c0c87ef6",
   430 => x"b7c08c4d",
   431 => x"87c603ac",
   432 => x"4da4c0c8",
   433 => x"efc24cc0",
   434 => x"49bf97e7",
   435 => x"d20299d0",
   436 => x"c21ec087",
   437 => x"fe49d6f5",
   438 => x"c487dec9",
   439 => x"4a497086",
   440 => x"c287efc0",
   441 => x"c21ef6e2",
   442 => x"fe49d6f5",
   443 => x"c487cac9",
   444 => x"4a497086",
   445 => x"c848d0ff",
   446 => x"d4c178c5",
   447 => x"bf976e7b",
   448 => x"c1486e7b",
   449 => x"c17e7080",
   450 => x"f0ff058d",
   451 => x"48d0ff87",
   452 => x"9a7278c4",
   453 => x"c087c505",
   454 => x"87e5c048",
   455 => x"f5c21ec1",
   456 => x"c6fe49d6",
   457 => x"86c487f2",
   458 => x"fe059c74",
   459 => x"d0ff87c4",
   460 => x"78c5c848",
   461 => x"c07bd3c1",
   462 => x"c178c47b",
   463 => x"c087c248",
   464 => x"4d262648",
   465 => x"4b264c26",
   466 => x"5e0e4f26",
   467 => x"710e5c5b",
   468 => x"0266cc4b",
   469 => x"4c87e8c0",
   470 => x"028cf0c0",
   471 => x"7487e8c0",
   472 => x"028ac14a",
   473 => x"8a87e0c0",
   474 => x"8a87dc02",
   475 => x"c087d802",
   476 => x"c0028ae0",
   477 => x"8ac187e3",
   478 => x"87e4c002",
   479 => x"7387e8c0",
   480 => x"87d9fb49",
   481 => x"7487e2c0",
   482 => x"f949c01e",
   483 => x"1e7487ca",
   484 => x"c3f94973",
   485 => x"d086c887",
   486 => x"c1497387",
   487 => x"87c987e9",
   488 => x"d5c24973",
   489 => x"c087c287",
   490 => x"87d8fe48",
   491 => x"e1c21e00",
   492 => x"c149bfef",
   493 => x"f3e1c2b9",
   494 => x"48d4ff59",
   495 => x"ff78ffc3",
   496 => x"e1c848d0",
   497 => x"48d4ff78",
   498 => x"31c478c1",
   499 => x"d0ff7871",
   500 => x"78e0c048",
   501 => x"711e4f26",
   502 => x"49a2c44a",
   503 => x"48ddf3c2",
   504 => x"4969786a",
   505 => x"e1c2b9c1",
   506 => x"c0ff59f3",
   507 => x"c6d0ff87",
   508 => x"2648c187",
   509 => x"4a711e4f",
   510 => x"c249a2c4",
   511 => x"7abfddf3",
   512 => x"bfefe1c2",
   513 => x"1e4f2679",
   514 => x"c21e4a71",
   515 => x"fe49d6f5",
   516 => x"c487cac1",
   517 => x"02987086",
   518 => x"e2c287dc",
   519 => x"f5c21ef6",
   520 => x"c4fe49d6",
   521 => x"86c487d3",
   522 => x"c9029870",
   523 => x"f6e2c287",
   524 => x"87e2fe49",
   525 => x"48c087c2",
   526 => x"711e4f26",
   527 => x"f5c21e4a",
   528 => x"c0fe49d6",
   529 => x"86c487d7",
   530 => x"de029870",
   531 => x"f6e2c287",
   532 => x"87e1fe49",
   533 => x"1ef6e2c2",
   534 => x"49d6f5c2",
   535 => x"87dcc4fe",
   536 => x"987086c4",
   537 => x"c187c402",
   538 => x"c087c248",
   539 => x"004f2648",
   540 => x"1e000000",
   541 => x"bfc0e2c2",
   542 => x"87e1f749",
   543 => x"4f2648c0",
   544 => x"00002884",
   545 => x"54534d41",
   546 => x"20444152",
   547 => x"004d4f52",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
