
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"48",x"d0",x"ff",x"1e"),
     1 => (x"71",x"78",x"e1",x"c8"),
     2 => (x"08",x"d4",x"ff",x"48"),
     3 => (x"1e",x"4f",x"26",x"78"),
     4 => (x"c8",x"48",x"d0",x"ff"),
     5 => (x"48",x"71",x"78",x"e1"),
     6 => (x"78",x"08",x"d4",x"ff"),
     7 => (x"ff",x"48",x"66",x"c4"),
     8 => (x"26",x"78",x"08",x"d4"),
     9 => (x"4a",x"71",x"1e",x"4f"),
    10 => (x"1e",x"49",x"66",x"c4"),
    11 => (x"de",x"ff",x"49",x"72"),
    12 => (x"48",x"d0",x"ff",x"87"),
    13 => (x"fc",x"78",x"e0",x"c0"),
    14 => (x"1e",x"4f",x"26",x"8e"),
    15 => (x"4a",x"71",x"1e",x"73"),
    16 => (x"ab",x"b7",x"c2",x"4b"),
    17 => (x"a3",x"87",x"c8",x"03"),
    18 => (x"ff",x"c3",x"4a",x"49"),
    19 => (x"ce",x"87",x"c7",x"9a"),
    20 => (x"c3",x"4a",x"49",x"a3"),
    21 => (x"66",x"c8",x"9a",x"ff"),
    22 => (x"49",x"72",x"1e",x"49"),
    23 => (x"fc",x"87",x"c6",x"ff"),
    24 => (x"26",x"4b",x"26",x"8e"),
    25 => (x"d0",x"ff",x"1e",x"4f"),
    26 => (x"78",x"c9",x"c8",x"48"),
    27 => (x"d4",x"ff",x"48",x"71"),
    28 => (x"4f",x"26",x"78",x"08"),
    29 => (x"49",x"4a",x"71",x"1e"),
    30 => (x"d0",x"ff",x"87",x"eb"),
    31 => (x"26",x"78",x"c8",x"48"),
    32 => (x"1e",x"73",x"1e",x"4f"),
    33 => (x"fc",x"c2",x"4b",x"71"),
    34 => (x"c3",x"02",x"bf",x"cc"),
    35 => (x"87",x"eb",x"c2",x"87"),
    36 => (x"c8",x"48",x"d0",x"ff"),
    37 => (x"48",x"73",x"78",x"c9"),
    38 => (x"ff",x"b0",x"e0",x"c0"),
    39 => (x"c2",x"78",x"08",x"d4"),
    40 => (x"c0",x"48",x"c0",x"fc"),
    41 => (x"02",x"66",x"c8",x"78"),
    42 => (x"ff",x"c3",x"87",x"c5"),
    43 => (x"c0",x"87",x"c2",x"49"),
    44 => (x"c8",x"fc",x"c2",x"49"),
    45 => (x"02",x"66",x"cc",x"59"),
    46 => (x"d5",x"c5",x"87",x"c6"),
    47 => (x"87",x"c4",x"4a",x"d5"),
    48 => (x"4a",x"ff",x"ff",x"cf"),
    49 => (x"5a",x"cc",x"fc",x"c2"),
    50 => (x"48",x"cc",x"fc",x"c2"),
    51 => (x"4b",x"26",x"78",x"c1"),
    52 => (x"5e",x"0e",x"4f",x"26"),
    53 => (x"0e",x"5d",x"5c",x"5b"),
    54 => (x"fc",x"c2",x"4d",x"71"),
    55 => (x"75",x"4b",x"bf",x"c8"),
    56 => (x"87",x"cb",x"02",x"9d"),
    57 => (x"c2",x"91",x"c8",x"49"),
    58 => (x"71",x"4a",x"f8",x"c1"),
    59 => (x"c2",x"87",x"c4",x"82"),
    60 => (x"c0",x"4a",x"f8",x"c5"),
    61 => (x"73",x"49",x"12",x"4c"),
    62 => (x"c4",x"fc",x"c2",x"99"),
    63 => (x"b8",x"71",x"48",x"bf"),
    64 => (x"78",x"08",x"d4",x"ff"),
    65 => (x"84",x"2b",x"b7",x"c1"),
    66 => (x"04",x"ac",x"b7",x"c8"),
    67 => (x"fc",x"c2",x"87",x"e7"),
    68 => (x"c8",x"48",x"bf",x"c0"),
    69 => (x"c4",x"fc",x"c2",x"80"),
    70 => (x"26",x"4d",x"26",x"58"),
    71 => (x"26",x"4b",x"26",x"4c"),
    72 => (x"1e",x"73",x"1e",x"4f"),
    73 => (x"4a",x"13",x"4b",x"71"),
    74 => (x"87",x"cb",x"02",x"9a"),
    75 => (x"e1",x"fe",x"49",x"72"),
    76 => (x"9a",x"4a",x"13",x"87"),
    77 => (x"26",x"87",x"f5",x"05"),
    78 => (x"1e",x"4f",x"26",x"4b"),
    79 => (x"bf",x"c0",x"fc",x"c2"),
    80 => (x"c0",x"fc",x"c2",x"49"),
    81 => (x"78",x"a1",x"c1",x"48"),
    82 => (x"a9",x"b7",x"c0",x"c4"),
    83 => (x"ff",x"87",x"db",x"03"),
    84 => (x"fc",x"c2",x"48",x"d4"),
    85 => (x"c2",x"78",x"bf",x"c4"),
    86 => (x"49",x"bf",x"c0",x"fc"),
    87 => (x"48",x"c0",x"fc",x"c2"),
    88 => (x"c4",x"78",x"a1",x"c1"),
    89 => (x"04",x"a9",x"b7",x"c0"),
    90 => (x"d0",x"ff",x"87",x"e5"),
    91 => (x"c2",x"78",x"c8",x"48"),
    92 => (x"c0",x"48",x"cc",x"fc"),
    93 => (x"00",x"4f",x"26",x"78"),
    94 => (x"00",x"00",x"00",x"00"),
    95 => (x"00",x"00",x"00",x"00"),
    96 => (x"5f",x"00",x"00",x"00"),
    97 => (x"00",x"00",x"00",x"5f"),
    98 => (x"00",x"03",x"03",x"00"),
    99 => (x"00",x"00",x"03",x"03"),
   100 => (x"14",x"7f",x"7f",x"14"),
   101 => (x"00",x"14",x"7f",x"7f"),
   102 => (x"6b",x"2e",x"24",x"00"),
   103 => (x"00",x"12",x"3a",x"6b"),
   104 => (x"18",x"36",x"6a",x"4c"),
   105 => (x"00",x"32",x"56",x"6c"),
   106 => (x"59",x"4f",x"7e",x"30"),
   107 => (x"40",x"68",x"3a",x"77"),
   108 => (x"07",x"04",x"00",x"00"),
   109 => (x"00",x"00",x"00",x"03"),
   110 => (x"3e",x"1c",x"00",x"00"),
   111 => (x"00",x"00",x"41",x"63"),
   112 => (x"63",x"41",x"00",x"00"),
   113 => (x"00",x"00",x"1c",x"3e"),
   114 => (x"1c",x"3e",x"2a",x"08"),
   115 => (x"08",x"2a",x"3e",x"1c"),
   116 => (x"3e",x"08",x"08",x"00"),
   117 => (x"00",x"08",x"08",x"3e"),
   118 => (x"e0",x"80",x"00",x"00"),
   119 => (x"00",x"00",x"00",x"60"),
   120 => (x"08",x"08",x"08",x"00"),
   121 => (x"00",x"08",x"08",x"08"),
   122 => (x"60",x"00",x"00",x"00"),
   123 => (x"00",x"00",x"00",x"60"),
   124 => (x"18",x"30",x"60",x"40"),
   125 => (x"01",x"03",x"06",x"0c"),
   126 => (x"59",x"7f",x"3e",x"00"),
   127 => (x"00",x"3e",x"7f",x"4d"),
   128 => (x"7f",x"06",x"04",x"00"),
   129 => (x"00",x"00",x"00",x"7f"),
   130 => (x"71",x"63",x"42",x"00"),
   131 => (x"00",x"46",x"4f",x"59"),
   132 => (x"49",x"63",x"22",x"00"),
   133 => (x"00",x"36",x"7f",x"49"),
   134 => (x"13",x"16",x"1c",x"18"),
   135 => (x"00",x"10",x"7f",x"7f"),
   136 => (x"45",x"67",x"27",x"00"),
   137 => (x"00",x"39",x"7d",x"45"),
   138 => (x"4b",x"7e",x"3c",x"00"),
   139 => (x"00",x"30",x"79",x"49"),
   140 => (x"71",x"01",x"01",x"00"),
   141 => (x"00",x"07",x"0f",x"79"),
   142 => (x"49",x"7f",x"36",x"00"),
   143 => (x"00",x"36",x"7f",x"49"),
   144 => (x"49",x"4f",x"06",x"00"),
   145 => (x"00",x"1e",x"3f",x"69"),
   146 => (x"66",x"00",x"00",x"00"),
   147 => (x"00",x"00",x"00",x"66"),
   148 => (x"e6",x"80",x"00",x"00"),
   149 => (x"00",x"00",x"00",x"66"),
   150 => (x"14",x"08",x"08",x"00"),
   151 => (x"00",x"22",x"22",x"14"),
   152 => (x"14",x"14",x"14",x"00"),
   153 => (x"00",x"14",x"14",x"14"),
   154 => (x"14",x"22",x"22",x"00"),
   155 => (x"00",x"08",x"08",x"14"),
   156 => (x"51",x"03",x"02",x"00"),
   157 => (x"00",x"06",x"0f",x"59"),
   158 => (x"5d",x"41",x"7f",x"3e"),
   159 => (x"00",x"1e",x"1f",x"55"),
   160 => (x"09",x"7f",x"7e",x"00"),
   161 => (x"00",x"7e",x"7f",x"09"),
   162 => (x"49",x"7f",x"7f",x"00"),
   163 => (x"00",x"36",x"7f",x"49"),
   164 => (x"63",x"3e",x"1c",x"00"),
   165 => (x"00",x"41",x"41",x"41"),
   166 => (x"41",x"7f",x"7f",x"00"),
   167 => (x"00",x"1c",x"3e",x"63"),
   168 => (x"49",x"7f",x"7f",x"00"),
   169 => (x"00",x"41",x"41",x"49"),
   170 => (x"09",x"7f",x"7f",x"00"),
   171 => (x"00",x"01",x"01",x"09"),
   172 => (x"41",x"7f",x"3e",x"00"),
   173 => (x"00",x"7a",x"7b",x"49"),
   174 => (x"08",x"7f",x"7f",x"00"),
   175 => (x"00",x"7f",x"7f",x"08"),
   176 => (x"7f",x"41",x"00",x"00"),
   177 => (x"00",x"00",x"41",x"7f"),
   178 => (x"40",x"60",x"20",x"00"),
   179 => (x"00",x"3f",x"7f",x"40"),
   180 => (x"1c",x"08",x"7f",x"7f"),
   181 => (x"00",x"41",x"63",x"36"),
   182 => (x"40",x"7f",x"7f",x"00"),
   183 => (x"00",x"40",x"40",x"40"),
   184 => (x"0c",x"06",x"7f",x"7f"),
   185 => (x"00",x"7f",x"7f",x"06"),
   186 => (x"0c",x"06",x"7f",x"7f"),
   187 => (x"00",x"7f",x"7f",x"18"),
   188 => (x"41",x"7f",x"3e",x"00"),
   189 => (x"00",x"3e",x"7f",x"41"),
   190 => (x"09",x"7f",x"7f",x"00"),
   191 => (x"00",x"06",x"0f",x"09"),
   192 => (x"61",x"41",x"7f",x"3e"),
   193 => (x"00",x"40",x"7e",x"7f"),
   194 => (x"09",x"7f",x"7f",x"00"),
   195 => (x"00",x"66",x"7f",x"19"),
   196 => (x"4d",x"6f",x"26",x"00"),
   197 => (x"00",x"32",x"7b",x"59"),
   198 => (x"7f",x"01",x"01",x"00"),
   199 => (x"00",x"01",x"01",x"7f"),
   200 => (x"40",x"7f",x"3f",x"00"),
   201 => (x"00",x"3f",x"7f",x"40"),
   202 => (x"70",x"3f",x"0f",x"00"),
   203 => (x"00",x"0f",x"3f",x"70"),
   204 => (x"18",x"30",x"7f",x"7f"),
   205 => (x"00",x"7f",x"7f",x"30"),
   206 => (x"1c",x"36",x"63",x"41"),
   207 => (x"41",x"63",x"36",x"1c"),
   208 => (x"7c",x"06",x"03",x"01"),
   209 => (x"01",x"03",x"06",x"7c"),
   210 => (x"4d",x"59",x"71",x"61"),
   211 => (x"00",x"41",x"43",x"47"),
   212 => (x"7f",x"7f",x"00",x"00"),
   213 => (x"00",x"00",x"41",x"41"),
   214 => (x"0c",x"06",x"03",x"01"),
   215 => (x"40",x"60",x"30",x"18"),
   216 => (x"41",x"41",x"00",x"00"),
   217 => (x"00",x"00",x"7f",x"7f"),
   218 => (x"03",x"06",x"0c",x"08"),
   219 => (x"00",x"08",x"0c",x"06"),
   220 => (x"80",x"80",x"80",x"80"),
   221 => (x"00",x"80",x"80",x"80"),
   222 => (x"03",x"00",x"00",x"00"),
   223 => (x"00",x"00",x"04",x"07"),
   224 => (x"54",x"74",x"20",x"00"),
   225 => (x"00",x"78",x"7c",x"54"),
   226 => (x"44",x"7f",x"7f",x"00"),
   227 => (x"00",x"38",x"7c",x"44"),
   228 => (x"44",x"7c",x"38",x"00"),
   229 => (x"00",x"00",x"44",x"44"),
   230 => (x"44",x"7c",x"38",x"00"),
   231 => (x"00",x"7f",x"7f",x"44"),
   232 => (x"54",x"7c",x"38",x"00"),
   233 => (x"00",x"18",x"5c",x"54"),
   234 => (x"7f",x"7e",x"04",x"00"),
   235 => (x"00",x"00",x"05",x"05"),
   236 => (x"a4",x"bc",x"18",x"00"),
   237 => (x"00",x"7c",x"fc",x"a4"),
   238 => (x"04",x"7f",x"7f",x"00"),
   239 => (x"00",x"78",x"7c",x"04"),
   240 => (x"3d",x"00",x"00",x"00"),
   241 => (x"00",x"00",x"40",x"7d"),
   242 => (x"80",x"80",x"80",x"00"),
   243 => (x"00",x"00",x"7d",x"fd"),
   244 => (x"10",x"7f",x"7f",x"00"),
   245 => (x"00",x"44",x"6c",x"38"),
   246 => (x"3f",x"00",x"00",x"00"),
   247 => (x"00",x"00",x"40",x"7f"),
   248 => (x"18",x"0c",x"7c",x"7c"),
   249 => (x"00",x"78",x"7c",x"0c"),
   250 => (x"04",x"7c",x"7c",x"00"),
   251 => (x"00",x"78",x"7c",x"04"),
   252 => (x"44",x"7c",x"38",x"00"),
   253 => (x"00",x"38",x"7c",x"44"),
   254 => (x"24",x"fc",x"fc",x"00"),
   255 => (x"00",x"18",x"3c",x"24"),
   256 => (x"24",x"3c",x"18",x"00"),
   257 => (x"00",x"fc",x"fc",x"24"),
   258 => (x"04",x"7c",x"7c",x"00"),
   259 => (x"00",x"08",x"0c",x"04"),
   260 => (x"54",x"5c",x"48",x"00"),
   261 => (x"00",x"20",x"74",x"54"),
   262 => (x"7f",x"3f",x"04",x"00"),
   263 => (x"00",x"00",x"44",x"44"),
   264 => (x"40",x"7c",x"3c",x"00"),
   265 => (x"00",x"7c",x"7c",x"40"),
   266 => (x"60",x"3c",x"1c",x"00"),
   267 => (x"00",x"1c",x"3c",x"60"),
   268 => (x"30",x"60",x"7c",x"3c"),
   269 => (x"00",x"3c",x"7c",x"60"),
   270 => (x"10",x"38",x"6c",x"44"),
   271 => (x"00",x"44",x"6c",x"38"),
   272 => (x"e0",x"bc",x"1c",x"00"),
   273 => (x"00",x"1c",x"3c",x"60"),
   274 => (x"74",x"64",x"44",x"00"),
   275 => (x"00",x"44",x"4c",x"5c"),
   276 => (x"3e",x"08",x"08",x"00"),
   277 => (x"00",x"41",x"41",x"77"),
   278 => (x"7f",x"00",x"00",x"00"),
   279 => (x"00",x"00",x"00",x"7f"),
   280 => (x"77",x"41",x"41",x"00"),
   281 => (x"00",x"08",x"08",x"3e"),
   282 => (x"03",x"01",x"01",x"02"),
   283 => (x"00",x"01",x"02",x"02"),
   284 => (x"7f",x"7f",x"7f",x"7f"),
   285 => (x"00",x"7f",x"7f",x"7f"),
   286 => (x"1c",x"1c",x"08",x"08"),
   287 => (x"7f",x"7f",x"3e",x"3e"),
   288 => (x"3e",x"3e",x"7f",x"7f"),
   289 => (x"08",x"08",x"1c",x"1c"),
   290 => (x"7c",x"18",x"10",x"00"),
   291 => (x"00",x"10",x"18",x"7c"),
   292 => (x"7c",x"30",x"10",x"00"),
   293 => (x"00",x"10",x"30",x"7c"),
   294 => (x"60",x"60",x"30",x"10"),
   295 => (x"00",x"06",x"1e",x"78"),
   296 => (x"18",x"3c",x"66",x"42"),
   297 => (x"00",x"42",x"66",x"3c"),
   298 => (x"c2",x"6a",x"38",x"78"),
   299 => (x"00",x"38",x"6c",x"c6"),
   300 => (x"60",x"00",x"00",x"60"),
   301 => (x"00",x"60",x"00",x"00"),
   302 => (x"5c",x"5b",x"5e",x"0e"),
   303 => (x"86",x"fc",x"0e",x"5d"),
   304 => (x"fc",x"c2",x"7e",x"71"),
   305 => (x"c0",x"4c",x"bf",x"d4"),
   306 => (x"c4",x"1e",x"c0",x"4b"),
   307 => (x"c4",x"02",x"ab",x"66"),
   308 => (x"c2",x"4d",x"c0",x"87"),
   309 => (x"75",x"4d",x"c1",x"87"),
   310 => (x"ee",x"49",x"73",x"1e"),
   311 => (x"86",x"c8",x"87",x"e3"),
   312 => (x"ef",x"49",x"e0",x"c0"),
   313 => (x"a4",x"c4",x"87",x"ec"),
   314 => (x"f0",x"49",x"6a",x"4a"),
   315 => (x"ca",x"f1",x"87",x"f3"),
   316 => (x"c1",x"84",x"cc",x"87"),
   317 => (x"ab",x"b7",x"c8",x"83"),
   318 => (x"87",x"cd",x"ff",x"04"),
   319 => (x"4d",x"26",x"8e",x"fc"),
   320 => (x"4b",x"26",x"4c",x"26"),
   321 => (x"71",x"1e",x"4f",x"26"),
   322 => (x"d8",x"fc",x"c2",x"4a"),
   323 => (x"d8",x"fc",x"c2",x"5a"),
   324 => (x"49",x"78",x"c7",x"48"),
   325 => (x"26",x"87",x"e1",x"fe"),
   326 => (x"1e",x"73",x"1e",x"4f"),
   327 => (x"b7",x"c0",x"4a",x"71"),
   328 => (x"87",x"d3",x"03",x"aa"),
   329 => (x"bf",x"fc",x"e0",x"c2"),
   330 => (x"c1",x"87",x"c4",x"05"),
   331 => (x"c0",x"87",x"c2",x"4b"),
   332 => (x"c0",x"e1",x"c2",x"4b"),
   333 => (x"c2",x"87",x"c4",x"5b"),
   334 => (x"fc",x"5a",x"c0",x"e1"),
   335 => (x"fc",x"e0",x"c2",x"48"),
   336 => (x"c1",x"4a",x"78",x"bf"),
   337 => (x"a2",x"c0",x"c1",x"9a"),
   338 => (x"87",x"e8",x"ec",x"49"),
   339 => (x"4f",x"26",x"4b",x"26"),
   340 => (x"c4",x"4a",x"71",x"1e"),
   341 => (x"49",x"72",x"1e",x"66"),
   342 => (x"fc",x"87",x"e0",x"eb"),
   343 => (x"1e",x"4f",x"26",x"8e"),
   344 => (x"c3",x"48",x"d4",x"ff"),
   345 => (x"d0",x"ff",x"78",x"ff"),
   346 => (x"78",x"e1",x"c0",x"48"),
   347 => (x"c1",x"48",x"d4",x"ff"),
   348 => (x"c4",x"48",x"71",x"78"),
   349 => (x"08",x"d4",x"ff",x"30"),
   350 => (x"48",x"d0",x"ff",x"78"),
   351 => (x"26",x"78",x"e0",x"c0"),
   352 => (x"5b",x"5e",x"0e",x"4f"),
   353 => (x"f0",x"0e",x"5d",x"5c"),
   354 => (x"48",x"a6",x"c8",x"86"),
   355 => (x"ec",x"4d",x"78",x"c0"),
   356 => (x"80",x"fc",x"7e",x"bf"),
   357 => (x"bf",x"d4",x"fc",x"c2"),
   358 => (x"4c",x"bf",x"e8",x"78"),
   359 => (x"bf",x"fc",x"e0",x"c2"),
   360 => (x"87",x"dd",x"e3",x"49"),
   361 => (x"ca",x"49",x"ee",x"cb"),
   362 => (x"4b",x"70",x"87",x"d6"),
   363 => (x"d2",x"e7",x"49",x"c7"),
   364 => (x"05",x"98",x"70",x"87"),
   365 => (x"49",x"6e",x"87",x"c8"),
   366 => (x"c1",x"02",x"99",x"c1"),
   367 => (x"4d",x"c1",x"87",x"c1"),
   368 => (x"c2",x"7e",x"bf",x"ec"),
   369 => (x"49",x"bf",x"fc",x"e0"),
   370 => (x"73",x"87",x"f6",x"e2"),
   371 => (x"87",x"fc",x"c9",x"49"),
   372 => (x"d7",x"02",x"98",x"70"),
   373 => (x"f4",x"e0",x"c2",x"87"),
   374 => (x"b9",x"c1",x"49",x"bf"),
   375 => (x"59",x"f8",x"e0",x"c2"),
   376 => (x"87",x"fb",x"fd",x"71"),
   377 => (x"c9",x"49",x"ee",x"cb"),
   378 => (x"4b",x"70",x"87",x"d6"),
   379 => (x"d2",x"e6",x"49",x"c7"),
   380 => (x"05",x"98",x"70",x"87"),
   381 => (x"6e",x"87",x"c7",x"ff"),
   382 => (x"05",x"99",x"c1",x"49"),
   383 => (x"75",x"87",x"ff",x"fe"),
   384 => (x"e3",x"c0",x"02",x"9d"),
   385 => (x"fc",x"e0",x"c2",x"87"),
   386 => (x"ba",x"c1",x"4a",x"bf"),
   387 => (x"5a",x"c0",x"e1",x"c2"),
   388 => (x"0a",x"7a",x"0a",x"fc"),
   389 => (x"c0",x"c1",x"9a",x"c1"),
   390 => (x"d7",x"e9",x"49",x"a2"),
   391 => (x"49",x"da",x"c1",x"87"),
   392 => (x"c8",x"87",x"e0",x"e5"),
   393 => (x"78",x"c1",x"48",x"a6"),
   394 => (x"bf",x"fc",x"e0",x"c2"),
   395 => (x"87",x"e9",x"c0",x"05"),
   396 => (x"ff",x"c3",x"49",x"74"),
   397 => (x"c0",x"1e",x"71",x"99"),
   398 => (x"87",x"d4",x"fc",x"49"),
   399 => (x"b7",x"c8",x"49",x"74"),
   400 => (x"c1",x"1e",x"71",x"29"),
   401 => (x"87",x"c8",x"fc",x"49"),
   402 => (x"fd",x"c3",x"86",x"c8"),
   403 => (x"87",x"f3",x"e4",x"49"),
   404 => (x"e4",x"49",x"fa",x"c3"),
   405 => (x"d1",x"c7",x"87",x"ed"),
   406 => (x"c3",x"49",x"74",x"87"),
   407 => (x"b7",x"c8",x"99",x"ff"),
   408 => (x"74",x"b4",x"71",x"2c"),
   409 => (x"87",x"df",x"02",x"9c"),
   410 => (x"bf",x"f8",x"e0",x"c2"),
   411 => (x"87",x"dc",x"c7",x"49"),
   412 => (x"c0",x"05",x"98",x"70"),
   413 => (x"4c",x"c0",x"87",x"c4"),
   414 => (x"e0",x"c2",x"87",x"d3"),
   415 => (x"87",x"c0",x"c7",x"49"),
   416 => (x"58",x"fc",x"e0",x"c2"),
   417 => (x"c2",x"87",x"c6",x"c0"),
   418 => (x"c0",x"48",x"f8",x"e0"),
   419 => (x"c8",x"49",x"74",x"78"),
   420 => (x"87",x"ce",x"05",x"99"),
   421 => (x"e3",x"49",x"f5",x"c3"),
   422 => (x"49",x"70",x"87",x"e9"),
   423 => (x"c0",x"02",x"99",x"c2"),
   424 => (x"fc",x"c2",x"87",x"e9"),
   425 => (x"c0",x"02",x"bf",x"d8"),
   426 => (x"c1",x"48",x"87",x"c9"),
   427 => (x"dc",x"fc",x"c2",x"88"),
   428 => (x"c4",x"87",x"d3",x"58"),
   429 => (x"e0",x"c1",x"48",x"66"),
   430 => (x"6e",x"7e",x"70",x"80"),
   431 => (x"c5",x"c0",x"02",x"bf"),
   432 => (x"49",x"ff",x"4b",x"87"),
   433 => (x"a6",x"c8",x"0f",x"73"),
   434 => (x"74",x"78",x"c1",x"48"),
   435 => (x"05",x"99",x"c4",x"49"),
   436 => (x"c3",x"87",x"ce",x"c0"),
   437 => (x"ea",x"e2",x"49",x"f2"),
   438 => (x"c2",x"49",x"70",x"87"),
   439 => (x"f0",x"c0",x"02",x"99"),
   440 => (x"d8",x"fc",x"c2",x"87"),
   441 => (x"c7",x"48",x"7e",x"bf"),
   442 => (x"c0",x"03",x"a8",x"b7"),
   443 => (x"48",x"6e",x"87",x"cb"),
   444 => (x"fc",x"c2",x"80",x"c1"),
   445 => (x"d3",x"c0",x"58",x"dc"),
   446 => (x"48",x"66",x"c4",x"87"),
   447 => (x"70",x"80",x"e0",x"c1"),
   448 => (x"02",x"bf",x"6e",x"7e"),
   449 => (x"4b",x"87",x"c5",x"c0"),
   450 => (x"0f",x"73",x"49",x"fe"),
   451 => (x"c1",x"48",x"a6",x"c8"),
   452 => (x"49",x"fd",x"c3",x"78"),
   453 => (x"70",x"87",x"ec",x"e1"),
   454 => (x"02",x"99",x"c2",x"49"),
   455 => (x"c2",x"87",x"e9",x"c0"),
   456 => (x"02",x"bf",x"d8",x"fc"),
   457 => (x"c2",x"87",x"c9",x"c0"),
   458 => (x"c0",x"48",x"d8",x"fc"),
   459 => (x"87",x"d3",x"c0",x"78"),
   460 => (x"c1",x"48",x"66",x"c4"),
   461 => (x"7e",x"70",x"80",x"e0"),
   462 => (x"c0",x"02",x"bf",x"6e"),
   463 => (x"fd",x"4b",x"87",x"c5"),
   464 => (x"c8",x"0f",x"73",x"49"),
   465 => (x"78",x"c1",x"48",x"a6"),
   466 => (x"e0",x"49",x"fa",x"c3"),
   467 => (x"49",x"70",x"87",x"f5"),
   468 => (x"c0",x"02",x"99",x"c2"),
   469 => (x"fc",x"c2",x"87",x"ea"),
   470 => (x"c7",x"48",x"bf",x"d8"),
   471 => (x"c0",x"03",x"a8",x"b7"),
   472 => (x"fc",x"c2",x"87",x"c9"),
   473 => (x"78",x"c7",x"48",x"d8"),
   474 => (x"c4",x"87",x"d0",x"c0"),
   475 => (x"e0",x"c1",x"4a",x"66"),
   476 => (x"c0",x"02",x"6a",x"82"),
   477 => (x"fc",x"4b",x"87",x"c5"),
   478 => (x"c8",x"0f",x"73",x"49"),
   479 => (x"78",x"c1",x"48",x"a6"),
   480 => (x"fc",x"c2",x"4d",x"c0"),
   481 => (x"50",x"c0",x"48",x"d0"),
   482 => (x"c2",x"49",x"ee",x"cb"),
   483 => (x"4b",x"70",x"87",x"f2"),
   484 => (x"97",x"d0",x"fc",x"c2"),
   485 => (x"dd",x"c1",x"05",x"bf"),
   486 => (x"c3",x"49",x"74",x"87"),
   487 => (x"c0",x"05",x"99",x"f0"),
   488 => (x"da",x"c1",x"87",x"cd"),
   489 => (x"da",x"df",x"ff",x"49"),
   490 => (x"02",x"98",x"70",x"87"),
   491 => (x"c1",x"87",x"c7",x"c1"),
   492 => (x"4c",x"bf",x"e8",x"4d"),
   493 => (x"99",x"ff",x"c3",x"49"),
   494 => (x"71",x"2c",x"b7",x"c8"),
   495 => (x"fc",x"e0",x"c2",x"b4"),
   496 => (x"da",x"ff",x"49",x"bf"),
   497 => (x"49",x"73",x"87",x"fb"),
   498 => (x"70",x"87",x"c1",x"c2"),
   499 => (x"c6",x"c0",x"02",x"98"),
   500 => (x"d0",x"fc",x"c2",x"87"),
   501 => (x"c2",x"50",x"c1",x"48"),
   502 => (x"bf",x"97",x"d0",x"fc"),
   503 => (x"87",x"d6",x"c0",x"05"),
   504 => (x"f0",x"c3",x"49",x"74"),
   505 => (x"c6",x"ff",x"05",x"99"),
   506 => (x"49",x"da",x"c1",x"87"),
   507 => (x"87",x"d3",x"de",x"ff"),
   508 => (x"fe",x"05",x"98",x"70"),
   509 => (x"9d",x"75",x"87",x"f9"),
   510 => (x"87",x"e0",x"c0",x"02"),
   511 => (x"c2",x"48",x"a6",x"cc"),
   512 => (x"78",x"bf",x"d8",x"fc"),
   513 => (x"cc",x"49",x"66",x"cc"),
   514 => (x"48",x"66",x"c4",x"91"),
   515 => (x"7e",x"70",x"80",x"71"),
   516 => (x"c0",x"02",x"bf",x"6e"),
   517 => (x"cc",x"4b",x"87",x"c6"),
   518 => (x"0f",x"73",x"49",x"66"),
   519 => (x"c0",x"02",x"66",x"c8"),
   520 => (x"fc",x"c2",x"87",x"c8"),
   521 => (x"f2",x"49",x"bf",x"d8"),
   522 => (x"8e",x"f0",x"87",x"ce"),
   523 => (x"4c",x"26",x"4d",x"26"),
   524 => (x"4f",x"26",x"4b",x"26"),
   525 => (x"00",x"00",x"00",x"00"),
   526 => (x"00",x"00",x"00",x"00"),
   527 => (x"00",x"00",x"00",x"00"),
   528 => (x"ff",x"4a",x"71",x"1e"),
   529 => (x"72",x"49",x"bf",x"c8"),
   530 => (x"4f",x"26",x"48",x"a1"),
   531 => (x"bf",x"c8",x"ff",x"1e"),
   532 => (x"c0",x"c0",x"fe",x"89"),
   533 => (x"a9",x"c0",x"c0",x"c0"),
   534 => (x"c0",x"87",x"c4",x"01"),
   535 => (x"c1",x"87",x"c2",x"4a"),
   536 => (x"26",x"48",x"72",x"4a"),
   537 => (x"5b",x"5e",x"0e",x"4f"),
   538 => (x"71",x"0e",x"5d",x"5c"),
   539 => (x"4c",x"d4",x"ff",x"4b"),
   540 => (x"c0",x"48",x"66",x"d0"),
   541 => (x"ff",x"49",x"d6",x"78"),
   542 => (x"c3",x"87",x"c5",x"de"),
   543 => (x"49",x"6c",x"7c",x"ff"),
   544 => (x"71",x"99",x"ff",x"c3"),
   545 => (x"f0",x"c3",x"49",x"4d"),
   546 => (x"a9",x"e0",x"c1",x"99"),
   547 => (x"c3",x"87",x"cb",x"05"),
   548 => (x"48",x"6c",x"7c",x"ff"),
   549 => (x"66",x"d0",x"98",x"c3"),
   550 => (x"ff",x"c3",x"78",x"08"),
   551 => (x"49",x"4a",x"6c",x"7c"),
   552 => (x"ff",x"c3",x"31",x"c8"),
   553 => (x"71",x"4a",x"6c",x"7c"),
   554 => (x"c8",x"49",x"72",x"b2"),
   555 => (x"7c",x"ff",x"c3",x"31"),
   556 => (x"b2",x"71",x"4a",x"6c"),
   557 => (x"31",x"c8",x"49",x"72"),
   558 => (x"6c",x"7c",x"ff",x"c3"),
   559 => (x"ff",x"b2",x"71",x"4a"),
   560 => (x"e0",x"c0",x"48",x"d0"),
   561 => (x"02",x"9b",x"73",x"78"),
   562 => (x"7b",x"72",x"87",x"c2"),
   563 => (x"4d",x"26",x"48",x"75"),
   564 => (x"4b",x"26",x"4c",x"26"),
   565 => (x"26",x"1e",x"4f",x"26"),
   566 => (x"5b",x"5e",x"0e",x"4f"),
   567 => (x"86",x"f8",x"0e",x"5c"),
   568 => (x"a6",x"c8",x"1e",x"76"),
   569 => (x"87",x"fd",x"fd",x"49"),
   570 => (x"4b",x"70",x"86",x"c4"),
   571 => (x"a8",x"c4",x"48",x"6e"),
   572 => (x"87",x"f4",x"c2",x"03"),
   573 => (x"f0",x"c3",x"4a",x"73"),
   574 => (x"aa",x"d0",x"c1",x"9a"),
   575 => (x"c1",x"87",x"c7",x"02"),
   576 => (x"c2",x"05",x"aa",x"e0"),
   577 => (x"49",x"73",x"87",x"e2"),
   578 => (x"c3",x"02",x"99",x"c8"),
   579 => (x"87",x"c6",x"ff",x"87"),
   580 => (x"9c",x"c3",x"4c",x"73"),
   581 => (x"c1",x"05",x"ac",x"c2"),
   582 => (x"66",x"c4",x"87",x"c4"),
   583 => (x"71",x"31",x"c9",x"49"),
   584 => (x"4a",x"66",x"c4",x"1e"),
   585 => (x"c2",x"92",x"c8",x"c1"),
   586 => (x"72",x"49",x"dc",x"fc"),
   587 => (x"c0",x"cc",x"fe",x"81"),
   588 => (x"ff",x"49",x"d8",x"87"),
   589 => (x"c8",x"87",x"c9",x"db"),
   590 => (x"ea",x"c2",x"1e",x"c0"),
   591 => (x"e1",x"fd",x"49",x"c0"),
   592 => (x"d0",x"ff",x"87",x"fa"),
   593 => (x"78",x"e0",x"c0",x"48"),
   594 => (x"1e",x"c0",x"ea",x"c2"),
   595 => (x"c1",x"4a",x"66",x"cc"),
   596 => (x"fc",x"c2",x"92",x"c8"),
   597 => (x"81",x"72",x"49",x"dc"),
   598 => (x"87",x"ca",x"c7",x"fe"),
   599 => (x"ac",x"c1",x"86",x"cc"),
   600 => (x"87",x"c4",x"c1",x"05"),
   601 => (x"c9",x"49",x"66",x"c4"),
   602 => (x"c4",x"1e",x"71",x"31"),
   603 => (x"c8",x"c1",x"4a",x"66"),
   604 => (x"dc",x"fc",x"c2",x"92"),
   605 => (x"fe",x"81",x"72",x"49"),
   606 => (x"c2",x"87",x"f6",x"ca"),
   607 => (x"c8",x"1e",x"c0",x"ea"),
   608 => (x"c8",x"c1",x"4a",x"66"),
   609 => (x"dc",x"fc",x"c2",x"92"),
   610 => (x"fe",x"81",x"72",x"49"),
   611 => (x"d7",x"87",x"c8",x"c5"),
   612 => (x"eb",x"d9",x"ff",x"49"),
   613 => (x"1e",x"c0",x"c8",x"87"),
   614 => (x"49",x"c0",x"ea",x"c2"),
   615 => (x"87",x"f9",x"df",x"fd"),
   616 => (x"d0",x"ff",x"86",x"cc"),
   617 => (x"78",x"e0",x"c0",x"48"),
   618 => (x"4c",x"26",x"8e",x"f8"),
   619 => (x"4f",x"26",x"4b",x"26"),
   620 => (x"5c",x"5b",x"5e",x"0e"),
   621 => (x"86",x"fc",x"0e",x"5d"),
   622 => (x"d4",x"ff",x"4d",x"71"),
   623 => (x"7e",x"66",x"d4",x"4c"),
   624 => (x"a8",x"b7",x"c3",x"48"),
   625 => (x"87",x"e3",x"c1",x"01"),
   626 => (x"66",x"c4",x"1e",x"75"),
   627 => (x"93",x"c8",x"c1",x"4b"),
   628 => (x"83",x"dc",x"fc",x"c2"),
   629 => (x"fd",x"fd",x"49",x"73"),
   630 => (x"a3",x"c8",x"87",x"ff"),
   631 => (x"ff",x"49",x"69",x"49"),
   632 => (x"e1",x"c8",x"48",x"d0"),
   633 => (x"71",x"7c",x"dd",x"78"),
   634 => (x"98",x"ff",x"c3",x"48"),
   635 => (x"4a",x"71",x"7c",x"70"),
   636 => (x"72",x"2a",x"b7",x"c8"),
   637 => (x"98",x"ff",x"c3",x"48"),
   638 => (x"4a",x"71",x"7c",x"70"),
   639 => (x"72",x"2a",x"b7",x"d0"),
   640 => (x"98",x"ff",x"c3",x"48"),
   641 => (x"48",x"71",x"7c",x"70"),
   642 => (x"70",x"28",x"b7",x"d8"),
   643 => (x"7c",x"7c",x"c0",x"7c"),
   644 => (x"7c",x"7c",x"7c",x"7c"),
   645 => (x"7c",x"7c",x"7c",x"7c"),
   646 => (x"d0",x"ff",x"7c",x"7c"),
   647 => (x"78",x"e0",x"c0",x"48"),
   648 => (x"dc",x"1e",x"66",x"c4"),
   649 => (x"fc",x"d7",x"ff",x"49"),
   650 => (x"fc",x"86",x"c8",x"87"),
   651 => (x"26",x"4d",x"26",x"8e"),
   652 => (x"26",x"4b",x"26",x"4c"),
   653 => (x"e9",x"c2",x"1e",x"4f"),
   654 => (x"fe",x"49",x"bf",x"c4"),
   655 => (x"c0",x"87",x"ef",x"dc"),
   656 => (x"00",x"4f",x"26",x"48"),
   657 => (x"00",x"00",x"2a",x"48"),
   658 => (x"54",x"53",x"4d",x"41"),
   659 => (x"20",x"44",x"41",x"52"),
   660 => (x"00",x"4d",x"4f",x"52"),
   661 => (x"00",x"00",x"1d",x"97"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

