library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"ecf5c287",
    12 => x"86c0c64e",
    13 => x"49ecf5c2",
    14 => x"48d0e2c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087cedf",
    19 => x"1e87fc98",
    20 => x"4a7186fc",
    21 => x"6949c0ff",
    22 => x"98c0c448",
    23 => x"026e7e70",
    24 => x"797287f5",
    25 => x"268efc48",
    26 => x"1e721e4f",
    27 => x"48121e73",
    28 => x"87ca0211",
    29 => x"98dfc34b",
    30 => x"0288739b",
    31 => x"4b2687f0",
    32 => x"4f264a26",
    33 => x"721e731e",
    34 => x"048bc11e",
    35 => x"481287ca",
    36 => x"87c40211",
    37 => x"87f10288",
    38 => x"4b264a26",
    39 => x"741e4f26",
    40 => x"721e731e",
    41 => x"048bc11e",
    42 => x"481287d0",
    43 => x"87ca0211",
    44 => x"98dfc34c",
    45 => x"0288749c",
    46 => x"4a2687eb",
    47 => x"4c264b26",
    48 => x"731e4f26",
    49 => x"a9738148",
    50 => x"1287c502",
    51 => x"87f60553",
    52 => x"c41e4f26",
    53 => x"48714a66",
    54 => x"fb055112",
    55 => x"1e4f2687",
    56 => x"114a66c4",
    57 => x"08d4ff48",
    58 => x"058ac178",
    59 => x"4f2687f5",
    60 => x"4a66c41e",
    61 => x"c348d4ff",
    62 => x"516878ff",
    63 => x"f3058ac1",
    64 => x"1e4f2687",
    65 => x"d4ff1e73",
    66 => x"7bffc34b",
    67 => x"ffc34a6b",
    68 => x"c8496b7b",
    69 => x"c3b17232",
    70 => x"4a6b7bff",
    71 => x"b27131c8",
    72 => x"6b7bffc3",
    73 => x"7232c849",
    74 => x"c44871b1",
    75 => x"264d2687",
    76 => x"264b264c",
    77 => x"5b5e0e4f",
    78 => x"710e5d5c",
    79 => x"4cd4ff4a",
    80 => x"ffc34972",
    81 => x"c27c7199",
    82 => x"05bfd0e2",
    83 => x"66d087c8",
    84 => x"d430c948",
    85 => x"66d058a6",
    86 => x"c329d849",
    87 => x"7c7199ff",
    88 => x"d04966d0",
    89 => x"99ffc329",
    90 => x"66d07c71",
    91 => x"c329c849",
    92 => x"7c7199ff",
    93 => x"c34966d0",
    94 => x"7c7199ff",
    95 => x"29d04972",
    96 => x"7199ffc3",
    97 => x"c94b6c7c",
    98 => x"c34dfff0",
    99 => x"d005abff",
   100 => x"7cffc387",
   101 => x"8dc14b6c",
   102 => x"c387c602",
   103 => x"f002abff",
   104 => x"fe487387",
   105 => x"c01e87c7",
   106 => x"48d4ff49",
   107 => x"c178ffc3",
   108 => x"b7c8c381",
   109 => x"87f104a9",
   110 => x"731e4f26",
   111 => x"c487e71e",
   112 => x"c04bdff8",
   113 => x"f0ffc01e",
   114 => x"fd49f7c1",
   115 => x"86c487e7",
   116 => x"c005a8c1",
   117 => x"d4ff87ea",
   118 => x"78ffc348",
   119 => x"c0c0c0c1",
   120 => x"c01ec0c0",
   121 => x"e9c1f0e1",
   122 => x"87c9fd49",
   123 => x"987086c4",
   124 => x"ff87ca05",
   125 => x"ffc348d4",
   126 => x"cb48c178",
   127 => x"87e6fe87",
   128 => x"fe058bc1",
   129 => x"48c087fd",
   130 => x"1e87e6fc",
   131 => x"d4ff1e73",
   132 => x"78ffc348",
   133 => x"1ec04bd3",
   134 => x"c1f0ffc0",
   135 => x"d4fc49c1",
   136 => x"7086c487",
   137 => x"87ca0598",
   138 => x"c348d4ff",
   139 => x"48c178ff",
   140 => x"f1fd87cb",
   141 => x"058bc187",
   142 => x"c087dbff",
   143 => x"87f1fb48",
   144 => x"5c5b5e0e",
   145 => x"4cd4ff0e",
   146 => x"c687dbfd",
   147 => x"e1c01eea",
   148 => x"49c8c1f0",
   149 => x"c487defb",
   150 => x"02a8c186",
   151 => x"eafe87c8",
   152 => x"c148c087",
   153 => x"dafa87e2",
   154 => x"cf497087",
   155 => x"c699ffff",
   156 => x"c802a9ea",
   157 => x"87d3fe87",
   158 => x"cbc148c0",
   159 => x"7cffc387",
   160 => x"fc4bf1c0",
   161 => x"987087f4",
   162 => x"87ebc002",
   163 => x"ffc01ec0",
   164 => x"49fac1f0",
   165 => x"c487defa",
   166 => x"05987086",
   167 => x"ffc387d9",
   168 => x"c3496c7c",
   169 => x"7c7c7cff",
   170 => x"99c0c17c",
   171 => x"c187c402",
   172 => x"c087d548",
   173 => x"c287d148",
   174 => x"87c405ab",
   175 => x"87c848c0",
   176 => x"fe058bc1",
   177 => x"48c087fd",
   178 => x"1e87e4f9",
   179 => x"e2c21e73",
   180 => x"78c148d0",
   181 => x"d0ff4bc7",
   182 => x"fb78c248",
   183 => x"d0ff87c8",
   184 => x"c078c348",
   185 => x"d0e5c01e",
   186 => x"f949c0c1",
   187 => x"86c487c7",
   188 => x"c105a8c1",
   189 => x"abc24b87",
   190 => x"c087c505",
   191 => x"87f9c048",
   192 => x"ff058bc1",
   193 => x"f7fc87d0",
   194 => x"d4e2c287",
   195 => x"05987058",
   196 => x"1ec187cd",
   197 => x"c1f0ffc0",
   198 => x"d8f849d0",
   199 => x"ff86c487",
   200 => x"ffc348d4",
   201 => x"87e0c478",
   202 => x"58d8e2c2",
   203 => x"c248d0ff",
   204 => x"48d4ff78",
   205 => x"c178ffc3",
   206 => x"87f5f748",
   207 => x"5c5b5e0e",
   208 => x"4a710e5d",
   209 => x"ff4dffc3",
   210 => x"7c754cd4",
   211 => x"c448d0ff",
   212 => x"7c7578c3",
   213 => x"ffc01e72",
   214 => x"49d8c1f0",
   215 => x"c487d6f7",
   216 => x"02987086",
   217 => x"48c087c5",
   218 => x"7587f0c0",
   219 => x"7cfec37c",
   220 => x"d41ec0c8",
   221 => x"e6f54966",
   222 => x"7586c487",
   223 => x"757c757c",
   224 => x"e0dad87c",
   225 => x"6c7c754b",
   226 => x"c5059949",
   227 => x"058bc187",
   228 => x"7c7587f3",
   229 => x"c248d0ff",
   230 => x"f648c178",
   231 => x"ff1e87cf",
   232 => x"d0ff4ad4",
   233 => x"78d1c448",
   234 => x"c17affc3",
   235 => x"87f80589",
   236 => x"731e4f26",
   237 => x"c54b711e",
   238 => x"4adfcdee",
   239 => x"c348d4ff",
   240 => x"486878ff",
   241 => x"02a8fec3",
   242 => x"8ac187c5",
   243 => x"7287ed05",
   244 => x"87c5059a",
   245 => x"eac048c0",
   246 => x"029b7387",
   247 => x"66c887cc",
   248 => x"f449731e",
   249 => x"86c487ca",
   250 => x"66c887c6",
   251 => x"87eefe49",
   252 => x"c348d4ff",
   253 => x"737878ff",
   254 => x"87c5059b",
   255 => x"d048d0ff",
   256 => x"f448c178",
   257 => x"731e87eb",
   258 => x"c04a711e",
   259 => x"48d4ff4b",
   260 => x"ff78ffc3",
   261 => x"c3c448d0",
   262 => x"48d4ff78",
   263 => x"7278ffc3",
   264 => x"f0ffc01e",
   265 => x"f449d1c1",
   266 => x"86c487cb",
   267 => x"cd059870",
   268 => x"1ec0c887",
   269 => x"fd4966cc",
   270 => x"86c487f8",
   271 => x"d0ff4b70",
   272 => x"7378c248",
   273 => x"87e9f348",
   274 => x"5c5b5e0e",
   275 => x"1ec00e5d",
   276 => x"c1f0ffc0",
   277 => x"dcf349c9",
   278 => x"c21ed287",
   279 => x"fd49d8e2",
   280 => x"86c887d0",
   281 => x"84c14cc0",
   282 => x"04acb7d2",
   283 => x"e2c287f8",
   284 => x"49bf97d8",
   285 => x"c199c0c3",
   286 => x"c005a9c0",
   287 => x"e2c287e7",
   288 => x"49bf97df",
   289 => x"e2c231d0",
   290 => x"4abf97e0",
   291 => x"b17232c8",
   292 => x"97e1e2c2",
   293 => x"71b14abf",
   294 => x"ffffcf4c",
   295 => x"84c19cff",
   296 => x"e7c134ca",
   297 => x"e1e2c287",
   298 => x"c149bf97",
   299 => x"c299c631",
   300 => x"bf97e2e2",
   301 => x"2ab7c74a",
   302 => x"e2c2b172",
   303 => x"4abf97dd",
   304 => x"c29dcf4d",
   305 => x"bf97dee2",
   306 => x"ca9ac34a",
   307 => x"dfe2c232",
   308 => x"c24bbf97",
   309 => x"c2b27333",
   310 => x"bf97e0e2",
   311 => x"9bc0c34b",
   312 => x"732bb7c6",
   313 => x"c181c2b2",
   314 => x"70307148",
   315 => x"7548c149",
   316 => x"724d7030",
   317 => x"7184c14c",
   318 => x"b7c0c894",
   319 => x"87cc06ad",
   320 => x"2db734c1",
   321 => x"adb7c0c8",
   322 => x"87f4ff01",
   323 => x"dcf04874",
   324 => x"5b5e0e87",
   325 => x"f80e5d5c",
   326 => x"feeac286",
   327 => x"c278c048",
   328 => x"c01ef6e2",
   329 => x"87defb49",
   330 => x"987086c4",
   331 => x"c087c505",
   332 => x"87cec948",
   333 => x"7ec14dc0",
   334 => x"bfdbf2c0",
   335 => x"ece3c249",
   336 => x"4bc8714a",
   337 => x"7087fdec",
   338 => x"87c20598",
   339 => x"f2c07ec0",
   340 => x"c249bfd7",
   341 => x"714ac8e4",
   342 => x"e7ec4bc8",
   343 => x"05987087",
   344 => x"7ec087c2",
   345 => x"fdc0026e",
   346 => x"fce9c287",
   347 => x"eac24dbf",
   348 => x"7ebf9ff4",
   349 => x"ead6c548",
   350 => x"87c705a8",
   351 => x"bffce9c2",
   352 => x"6e87ce4d",
   353 => x"d5e9ca48",
   354 => x"87c502a8",
   355 => x"f1c748c0",
   356 => x"f6e2c287",
   357 => x"f949751e",
   358 => x"86c487ec",
   359 => x"c5059870",
   360 => x"c748c087",
   361 => x"f2c087dc",
   362 => x"c249bfd7",
   363 => x"714ac8e4",
   364 => x"cfeb4bc8",
   365 => x"05987087",
   366 => x"eac287c8",
   367 => x"78c148fe",
   368 => x"f2c087da",
   369 => x"c249bfdb",
   370 => x"714aece3",
   371 => x"f3ea4bc8",
   372 => x"02987087",
   373 => x"c087c5c0",
   374 => x"87e6c648",
   375 => x"97f4eac2",
   376 => x"d5c149bf",
   377 => x"cdc005a9",
   378 => x"f5eac287",
   379 => x"c249bf97",
   380 => x"c002a9ea",
   381 => x"48c087c5",
   382 => x"c287c7c6",
   383 => x"bf97f6e2",
   384 => x"e9c3487e",
   385 => x"cec002a8",
   386 => x"c3486e87",
   387 => x"c002a8eb",
   388 => x"48c087c5",
   389 => x"c287ebc5",
   390 => x"bf97c1e3",
   391 => x"c0059949",
   392 => x"e3c287cc",
   393 => x"49bf97c2",
   394 => x"c002a9c2",
   395 => x"48c087c5",
   396 => x"c287cfc5",
   397 => x"bf97c3e3",
   398 => x"faeac248",
   399 => x"484c7058",
   400 => x"eac288c1",
   401 => x"e3c258fe",
   402 => x"49bf97c4",
   403 => x"e3c28175",
   404 => x"4abf97c5",
   405 => x"a17232c8",
   406 => x"cbefc27e",
   407 => x"c2786e48",
   408 => x"bf97c6e3",
   409 => x"58a6c848",
   410 => x"bffeeac2",
   411 => x"87d4c202",
   412 => x"bfd7f2c0",
   413 => x"c8e4c249",
   414 => x"4bc8714a",
   415 => x"7087c5e8",
   416 => x"c5c00298",
   417 => x"c348c087",
   418 => x"eac287f8",
   419 => x"c24cbff6",
   420 => x"c25cdfef",
   421 => x"bf97dbe3",
   422 => x"c231c849",
   423 => x"bf97dae3",
   424 => x"c249a14a",
   425 => x"bf97dce3",
   426 => x"7232d04a",
   427 => x"e3c249a1",
   428 => x"4abf97dd",
   429 => x"a17232d8",
   430 => x"9166c449",
   431 => x"bfcbefc2",
   432 => x"d3efc281",
   433 => x"e3e3c259",
   434 => x"c84abf97",
   435 => x"e2e3c232",
   436 => x"a24bbf97",
   437 => x"e4e3c24a",
   438 => x"d04bbf97",
   439 => x"4aa27333",
   440 => x"97e5e3c2",
   441 => x"9bcf4bbf",
   442 => x"a27333d8",
   443 => x"d7efc24a",
   444 => x"d3efc25a",
   445 => x"8ac24abf",
   446 => x"efc29274",
   447 => x"a17248d7",
   448 => x"87cac178",
   449 => x"97c8e3c2",
   450 => x"31c849bf",
   451 => x"97c7e3c2",
   452 => x"49a14abf",
   453 => x"59c6ebc2",
   454 => x"bfc2ebc2",
   455 => x"c731c549",
   456 => x"29c981ff",
   457 => x"59dfefc2",
   458 => x"97cde3c2",
   459 => x"32c84abf",
   460 => x"97cce3c2",
   461 => x"4aa24bbf",
   462 => x"6e9266c4",
   463 => x"dbefc282",
   464 => x"d3efc25a",
   465 => x"c278c048",
   466 => x"7248cfef",
   467 => x"efc278a1",
   468 => x"efc248df",
   469 => x"c278bfd3",
   470 => x"c248e3ef",
   471 => x"78bfd7ef",
   472 => x"bffeeac2",
   473 => x"87c9c002",
   474 => x"30c44874",
   475 => x"c9c07e70",
   476 => x"dbefc287",
   477 => x"30c448bf",
   478 => x"ebc27e70",
   479 => x"786e48c2",
   480 => x"8ef848c1",
   481 => x"4c264d26",
   482 => x"4f264b26",
   483 => x"5c5b5e0e",
   484 => x"4a710e5d",
   485 => x"bffeeac2",
   486 => x"7287cb02",
   487 => x"722bc74b",
   488 => x"9cffc14c",
   489 => x"4b7287c9",
   490 => x"4c722bc8",
   491 => x"c29cffc3",
   492 => x"83bfcbef",
   493 => x"bfd3f2c0",
   494 => x"87d902ab",
   495 => x"5bd7f2c0",
   496 => x"1ef6e2c2",
   497 => x"fdf04973",
   498 => x"7086c487",
   499 => x"87c50598",
   500 => x"e6c048c0",
   501 => x"feeac287",
   502 => x"87d202bf",
   503 => x"91c44974",
   504 => x"81f6e2c2",
   505 => x"ffcf4d69",
   506 => x"9dffffff",
   507 => x"497487cb",
   508 => x"e2c291c2",
   509 => x"699f81f6",
   510 => x"fe48754d",
   511 => x"5e0e87c6",
   512 => x"0e5d5c5b",
   513 => x"c04d711e",
   514 => x"ca49c11e",
   515 => x"86c487ee",
   516 => x"029c4c70",
   517 => x"c287c0c1",
   518 => x"754ac6eb",
   519 => x"87c9e149",
   520 => x"c0029870",
   521 => x"4a7487f1",
   522 => x"4bcb4975",
   523 => x"7087efe1",
   524 => x"e2c00298",
   525 => x"741ec087",
   526 => x"87c7029c",
   527 => x"c048a6c4",
   528 => x"c487c578",
   529 => x"78c148a6",
   530 => x"c94966c4",
   531 => x"86c487ee",
   532 => x"059c4c70",
   533 => x"7487c0ff",
   534 => x"e7fc2648",
   535 => x"5b5e0e87",
   536 => x"1e0e5d5c",
   537 => x"059b4b71",
   538 => x"48c087c5",
   539 => x"c887e5c1",
   540 => x"7dc04da3",
   541 => x"c70266d4",
   542 => x"9766d487",
   543 => x"87c505bf",
   544 => x"cfc148c0",
   545 => x"4966d487",
   546 => x"7087f3fd",
   547 => x"c1029c4c",
   548 => x"a4dc87c0",
   549 => x"da7d6949",
   550 => x"a3c449a4",
   551 => x"7a699f4a",
   552 => x"bffeeac2",
   553 => x"d487d202",
   554 => x"699f49a4",
   555 => x"ffffc049",
   556 => x"d0487199",
   557 => x"c27e7030",
   558 => x"6e7ec087",
   559 => x"806a4849",
   560 => x"7bc07a70",
   561 => x"6a49a3cc",
   562 => x"49a3d079",
   563 => x"487479c0",
   564 => x"48c087c2",
   565 => x"87ecfa26",
   566 => x"5c5b5e0e",
   567 => x"4c710e5d",
   568 => x"48d3f2c0",
   569 => x"9c7478ff",
   570 => x"87cac102",
   571 => x"6949a4c8",
   572 => x"87c2c102",
   573 => x"6c4a66d0",
   574 => x"a6d48249",
   575 => x"4d66d05a",
   576 => x"faeac2b9",
   577 => x"baff4abf",
   578 => x"99719972",
   579 => x"87e4c002",
   580 => x"6b4ba4c4",
   581 => x"87f4f949",
   582 => x"eac27b70",
   583 => x"6c49bff6",
   584 => x"757c7181",
   585 => x"faeac2b9",
   586 => x"baff4abf",
   587 => x"99719972",
   588 => x"87dcff05",
   589 => x"cbf97c75",
   590 => x"1e731e87",
   591 => x"029b4b71",
   592 => x"a3c887c7",
   593 => x"c5056949",
   594 => x"c048c087",
   595 => x"efc287eb",
   596 => x"c44abfcf",
   597 => x"496949a3",
   598 => x"eac289c2",
   599 => x"7191bff6",
   600 => x"eac24aa2",
   601 => x"6b49bffa",
   602 => x"4aa27199",
   603 => x"721e66c8",
   604 => x"87d2ea49",
   605 => x"497086c4",
   606 => x"87ccf848",
   607 => x"711e731e",
   608 => x"c7029b4b",
   609 => x"49a3c887",
   610 => x"87c50569",
   611 => x"ebc048c0",
   612 => x"cfefc287",
   613 => x"a3c44abf",
   614 => x"c2496949",
   615 => x"f6eac289",
   616 => x"a27191bf",
   617 => x"faeac24a",
   618 => x"996b49bf",
   619 => x"c84aa271",
   620 => x"49721e66",
   621 => x"c487c5e6",
   622 => x"48497086",
   623 => x"0e87c9f7",
   624 => x"5d5c5b5e",
   625 => x"4b711e0e",
   626 => x"c94c66d4",
   627 => x"029b732c",
   628 => x"c887cfc1",
   629 => x"026949a3",
   630 => x"d087c7c1",
   631 => x"66d44da3",
   632 => x"faeac27d",
   633 => x"b9ff49bf",
   634 => x"7e994a6b",
   635 => x"cd03ac71",
   636 => x"7d7bc087",
   637 => x"c44aa3cc",
   638 => x"796a49a3",
   639 => x"8c7287c2",
   640 => x"dd029c74",
   641 => x"731e4987",
   642 => x"87ccfb49",
   643 => x"66d486c4",
   644 => x"99ffc749",
   645 => x"c287cb02",
   646 => x"731ef6e2",
   647 => x"87d9fc49",
   648 => x"f52686c4",
   649 => x"731e87de",
   650 => x"9b4b711e",
   651 => x"87e4c002",
   652 => x"5be3efc2",
   653 => x"8ac24a73",
   654 => x"bff6eac2",
   655 => x"efc29249",
   656 => x"7248bfcf",
   657 => x"e7efc280",
   658 => x"c4487158",
   659 => x"c6ebc230",
   660 => x"87edc058",
   661 => x"48dfefc2",
   662 => x"bfd3efc2",
   663 => x"e3efc278",
   664 => x"d7efc248",
   665 => x"eac278bf",
   666 => x"c902bffe",
   667 => x"f6eac287",
   668 => x"31c449bf",
   669 => x"efc287c7",
   670 => x"c449bfdb",
   671 => x"c6ebc231",
   672 => x"87c4f459",
   673 => x"5c5b5e0e",
   674 => x"c04a710e",
   675 => x"029a724b",
   676 => x"da87e1c0",
   677 => x"699f49a2",
   678 => x"feeac24b",
   679 => x"87cf02bf",
   680 => x"9f49a2d4",
   681 => x"c04c4969",
   682 => x"d09cffff",
   683 => x"c087c234",
   684 => x"b349744c",
   685 => x"edfd4973",
   686 => x"87caf387",
   687 => x"5c5b5e0e",
   688 => x"86f40e5d",
   689 => x"7ec04a71",
   690 => x"d8029a72",
   691 => x"f2e2c287",
   692 => x"c278c048",
   693 => x"c248eae2",
   694 => x"78bfe3ef",
   695 => x"48eee2c2",
   696 => x"bfdfefc2",
   697 => x"d3ebc278",
   698 => x"c250c048",
   699 => x"49bfc2eb",
   700 => x"bff2e2c2",
   701 => x"03aa714a",
   702 => x"7287ffc3",
   703 => x"0599cf49",
   704 => x"c287e0c0",
   705 => x"c21ef6e2",
   706 => x"49bfeae2",
   707 => x"48eae2c2",
   708 => x"7178a1c1",
   709 => x"c487efe3",
   710 => x"cff2c086",
   711 => x"f6e2c248",
   712 => x"c087cc78",
   713 => x"48bfcff2",
   714 => x"c080e0c0",
   715 => x"c258d3f2",
   716 => x"48bff2e2",
   717 => x"e2c280c1",
   718 => x"8f2758f6",
   719 => x"bf00000c",
   720 => x"9d4dbf97",
   721 => x"87e2c202",
   722 => x"02ade5c3",
   723 => x"c087dbc2",
   724 => x"4bbfcff2",
   725 => x"1149a3cb",
   726 => x"05accf4c",
   727 => x"7587d2c1",
   728 => x"c199df49",
   729 => x"c291cd89",
   730 => x"c181c6eb",
   731 => x"51124aa3",
   732 => x"124aa3c3",
   733 => x"4aa3c551",
   734 => x"a3c75112",
   735 => x"c951124a",
   736 => x"51124aa3",
   737 => x"124aa3ce",
   738 => x"4aa3d051",
   739 => x"a3d25112",
   740 => x"d451124a",
   741 => x"51124aa3",
   742 => x"124aa3d6",
   743 => x"4aa3d851",
   744 => x"a3dc5112",
   745 => x"de51124a",
   746 => x"51124aa3",
   747 => x"f9c07ec1",
   748 => x"c8497487",
   749 => x"eac00599",
   750 => x"d0497487",
   751 => x"87d00599",
   752 => x"c00266dc",
   753 => x"497387ca",
   754 => x"700f66dc",
   755 => x"87d30298",
   756 => x"c6c0056e",
   757 => x"c6ebc287",
   758 => x"c050c048",
   759 => x"48bfcff2",
   760 => x"c287e7c2",
   761 => x"c048d3eb",
   762 => x"ebc27e50",
   763 => x"c249bfc2",
   764 => x"4abff2e2",
   765 => x"fc04aa71",
   766 => x"efc287c1",
   767 => x"c005bfe3",
   768 => x"eac287c8",
   769 => x"c102bffe",
   770 => x"f2c087fe",
   771 => x"78ff48d3",
   772 => x"bfeee2c2",
   773 => x"87f4ed49",
   774 => x"e2c24970",
   775 => x"a6c459f2",
   776 => x"eee2c248",
   777 => x"eac278bf",
   778 => x"c002bffe",
   779 => x"66c487d8",
   780 => x"ffffcf49",
   781 => x"a999f8ff",
   782 => x"87c5c002",
   783 => x"e1c04dc0",
   784 => x"c04dc187",
   785 => x"66c487dc",
   786 => x"f8ffcf49",
   787 => x"c002a999",
   788 => x"a6c887c8",
   789 => x"c078c048",
   790 => x"a6c887c5",
   791 => x"c878c148",
   792 => x"9d754d66",
   793 => x"87e0c005",
   794 => x"c24966c4",
   795 => x"f6eac289",
   796 => x"c2914abf",
   797 => x"4abfcfef",
   798 => x"48eae2c2",
   799 => x"c278a172",
   800 => x"c048f2e2",
   801 => x"87e3f978",
   802 => x"8ef448c0",
   803 => x"0087f5eb",
   804 => x"ff000000",
   805 => x"9fffffff",
   806 => x"a800000c",
   807 => x"4600000c",
   808 => x"32335441",
   809 => x"00202020",
   810 => x"31544146",
   811 => x"20202036",
   812 => x"d4ff1e00",
   813 => x"78ffc348",
   814 => x"4f264868",
   815 => x"48d4ff1e",
   816 => x"ff78ffc3",
   817 => x"e1c848d0",
   818 => x"48d4ff78",
   819 => x"efc278d4",
   820 => x"d4ff48e7",
   821 => x"4f2650bf",
   822 => x"48d0ff1e",
   823 => x"2678e0c0",
   824 => x"ccff1e4f",
   825 => x"99497087",
   826 => x"c087c602",
   827 => x"f105a9fb",
   828 => x"26487187",
   829 => x"5b5e0e4f",
   830 => x"4b710e5c",
   831 => x"f0fe4cc0",
   832 => x"99497087",
   833 => x"87f9c002",
   834 => x"02a9ecc0",
   835 => x"c087f2c0",
   836 => x"c002a9fb",
   837 => x"66cc87eb",
   838 => x"c703acb7",
   839 => x"0266d087",
   840 => x"537187c2",
   841 => x"c2029971",
   842 => x"fe84c187",
   843 => x"497087c3",
   844 => x"87cd0299",
   845 => x"02a9ecc0",
   846 => x"fbc087c7",
   847 => x"d5ff05a9",
   848 => x"0266d087",
   849 => x"97c087c3",
   850 => x"a9ecc07b",
   851 => x"7487c405",
   852 => x"7487c54a",
   853 => x"8a0ac04a",
   854 => x"87c24872",
   855 => x"4c264d26",
   856 => x"4f264b26",
   857 => x"87c9fd1e",
   858 => x"f0c04970",
   859 => x"ca04a9b7",
   860 => x"b7f9c087",
   861 => x"87c301a9",
   862 => x"c189f0c0",
   863 => x"04a9b7c1",
   864 => x"dac187ca",
   865 => x"c301a9b7",
   866 => x"89f7c087",
   867 => x"4f264871",
   868 => x"5c5b5e0e",
   869 => x"ff4a710e",
   870 => x"49724cd4",
   871 => x"7087eac0",
   872 => x"c2029b4b",
   873 => x"ff8bc187",
   874 => x"c5c848d0",
   875 => x"7cd5c178",
   876 => x"31c64973",
   877 => x"97ecdec2",
   878 => x"71484abf",
   879 => x"ff7c70b0",
   880 => x"78c448d0",
   881 => x"d5fe4873",
   882 => x"5b5e0e87",
   883 => x"f80e5d5c",
   884 => x"c04b7186",
   885 => x"f0fac07e",
   886 => x"df49bf97",
   887 => x"eec005a9",
   888 => x"49a3c887",
   889 => x"c1496997",
   890 => x"dd05a9c3",
   891 => x"49a3c987",
   892 => x"c1496997",
   893 => x"d105a9c6",
   894 => x"49a3ca87",
   895 => x"c1496997",
   896 => x"c505a9c7",
   897 => x"c248c187",
   898 => x"48c087e1",
   899 => x"fa87dcc2",
   900 => x"4cc087ea",
   901 => x"97f0fac0",
   902 => x"a9c049bf",
   903 => x"fa87cf04",
   904 => x"84c187ff",
   905 => x"97f0fac0",
   906 => x"06ac49bf",
   907 => x"fac087f1",
   908 => x"02bf97f0",
   909 => x"f8f987cf",
   910 => x"99497087",
   911 => x"c087c602",
   912 => x"f105a9ec",
   913 => x"f94cc087",
   914 => x"4d7087e7",
   915 => x"c887e2f9",
   916 => x"dcf958a6",
   917 => x"c14a7087",
   918 => x"49a3c884",
   919 => x"ad496997",
   920 => x"c087c702",
   921 => x"c005adff",
   922 => x"a3c987e7",
   923 => x"49699749",
   924 => x"02a966c4",
   925 => x"c04887c7",
   926 => x"d405a8ff",
   927 => x"49a3ca87",
   928 => x"aa496997",
   929 => x"c087c602",
   930 => x"c405aaff",
   931 => x"d07ec187",
   932 => x"adecc087",
   933 => x"c087c602",
   934 => x"c405adfb",
   935 => x"c14cc087",
   936 => x"fe026e7e",
   937 => x"eff887e1",
   938 => x"f8487487",
   939 => x"87ecfa8e",
   940 => x"5b5e0e00",
   941 => x"1e0e5d5c",
   942 => x"4cc04b71",
   943 => x"c004ab4d",
   944 => x"f7c087e8",
   945 => x"9d751ec9",
   946 => x"c087c402",
   947 => x"c187c24a",
   948 => x"ef49724a",
   949 => x"86c487e6",
   950 => x"84c17e70",
   951 => x"87c2056e",
   952 => x"85c14c73",
   953 => x"ff06ac73",
   954 => x"486e87d8",
   955 => x"264d2626",
   956 => x"264b264c",
   957 => x"5b5e0e4f",
   958 => x"1e0e5d5c",
   959 => x"de494c71",
   960 => x"c1f0c291",
   961 => x"9785714d",
   962 => x"ddc1026d",
   963 => x"ecefc287",
   964 => x"82744abf",
   965 => x"d8fe4972",
   966 => x"6e7e7087",
   967 => x"87f3c002",
   968 => x"4bf4efc2",
   969 => x"49cb4a6e",
   970 => x"87d6c6ff",
   971 => x"93cb4b74",
   972 => x"83e0e1c1",
   973 => x"fdc083c4",
   974 => x"49747bee",
   975 => x"87f7c5c1",
   976 => x"f0c27b75",
   977 => x"49bf97c0",
   978 => x"f4efc21e",
   979 => x"f9dfc149",
   980 => x"7486c487",
   981 => x"dec5c149",
   982 => x"c149c087",
   983 => x"c287fdc6",
   984 => x"c048e8ef",
   985 => x"df49c178",
   986 => x"fd2687fd",
   987 => x"6f4c87ff",
   988 => x"6e696461",
   989 => x"2e2e2e67",
   990 => x"5b5e0e00",
   991 => x"4b710e5c",
   992 => x"ecefc24a",
   993 => x"497282bf",
   994 => x"7087e6fc",
   995 => x"c4029c4c",
   996 => x"efeb4987",
   997 => x"ecefc287",
   998 => x"c178c048",
   999 => x"87c7df49",
  1000 => x"0e87ccfd",
  1001 => x"5d5c5b5e",
  1002 => x"c286f40e",
  1003 => x"c04df6e2",
  1004 => x"48a6c44c",
  1005 => x"efc278c0",
  1006 => x"c049bfec",
  1007 => x"c1c106a9",
  1008 => x"f6e2c287",
  1009 => x"c0029848",
  1010 => x"f7c087f8",
  1011 => x"66c81ec9",
  1012 => x"c487c702",
  1013 => x"78c048a6",
  1014 => x"a6c487c5",
  1015 => x"c478c148",
  1016 => x"d7eb4966",
  1017 => x"7086c487",
  1018 => x"c484c14d",
  1019 => x"80c14866",
  1020 => x"c258a6c8",
  1021 => x"49bfecef",
  1022 => x"87c603ac",
  1023 => x"ff059d75",
  1024 => x"4cc087c8",
  1025 => x"c3029d75",
  1026 => x"f7c087e0",
  1027 => x"66c81ec9",
  1028 => x"cc87c702",
  1029 => x"78c048a6",
  1030 => x"a6cc87c5",
  1031 => x"cc78c148",
  1032 => x"d7ea4966",
  1033 => x"7086c487",
  1034 => x"c2026e7e",
  1035 => x"496e87e9",
  1036 => x"699781cb",
  1037 => x"0299d049",
  1038 => x"c087d6c1",
  1039 => x"744af9fd",
  1040 => x"c191cb49",
  1041 => x"7281e0e1",
  1042 => x"c381c879",
  1043 => x"497451ff",
  1044 => x"f0c291de",
  1045 => x"85714dc1",
  1046 => x"7d97c1c2",
  1047 => x"c049a5c1",
  1048 => x"ebc251e0",
  1049 => x"02bf97c6",
  1050 => x"84c187d2",
  1051 => x"c24ba5c2",
  1052 => x"db4ac6eb",
  1053 => x"c9c1ff49",
  1054 => x"87dbc187",
  1055 => x"c049a5cd",
  1056 => x"c284c151",
  1057 => x"4a6e4ba5",
  1058 => x"c0ff49cb",
  1059 => x"c6c187f4",
  1060 => x"f5fbc087",
  1061 => x"cb49744a",
  1062 => x"e0e1c191",
  1063 => x"c2797281",
  1064 => x"bf97c6eb",
  1065 => x"7487d802",
  1066 => x"c191de49",
  1067 => x"c1f0c284",
  1068 => x"c283714b",
  1069 => x"dd4ac6eb",
  1070 => x"c5c0ff49",
  1071 => x"7487d887",
  1072 => x"c293de4b",
  1073 => x"cb83c1f0",
  1074 => x"51c049a3",
  1075 => x"6e7384c1",
  1076 => x"fe49cb4a",
  1077 => x"c487ebff",
  1078 => x"80c14866",
  1079 => x"c758a6c8",
  1080 => x"c5c003ac",
  1081 => x"fc056e87",
  1082 => x"487487e0",
  1083 => x"fcf78ef4",
  1084 => x"1e731e87",
  1085 => x"cb494b71",
  1086 => x"e0e1c191",
  1087 => x"4aa1c881",
  1088 => x"48ecdec2",
  1089 => x"a1c95012",
  1090 => x"f0fac04a",
  1091 => x"ca501248",
  1092 => x"c0f0c281",
  1093 => x"c2501148",
  1094 => x"bf97c0f0",
  1095 => x"49c01e49",
  1096 => x"87e6d8c1",
  1097 => x"48e8efc2",
  1098 => x"49c178de",
  1099 => x"2687f8d8",
  1100 => x"1e87fef6",
  1101 => x"cb494a71",
  1102 => x"e0e1c191",
  1103 => x"1181c881",
  1104 => x"ecefc248",
  1105 => x"ecefc258",
  1106 => x"c178c048",
  1107 => x"87d7d849",
  1108 => x"c01e4f26",
  1109 => x"c3ffc049",
  1110 => x"1e4f2687",
  1111 => x"d2029971",
  1112 => x"f5e2c187",
  1113 => x"f750c048",
  1114 => x"f3c4c180",
  1115 => x"cee1c140",
  1116 => x"c187ce78",
  1117 => x"c148f1e2",
  1118 => x"fc78efe0",
  1119 => x"d2c5c180",
  1120 => x"0e4f2678",
  1121 => x"0e5c5b5e",
  1122 => x"cb4a4c71",
  1123 => x"e0e1c192",
  1124 => x"49a2c882",
  1125 => x"974ba2c9",
  1126 => x"971e4b6b",
  1127 => x"ca1e4969",
  1128 => x"c0491282",
  1129 => x"c087fee9",
  1130 => x"87fbd649",
  1131 => x"fcc04974",
  1132 => x"8ef887c5",
  1133 => x"1e87f8f4",
  1134 => x"4b711e73",
  1135 => x"87c3ff49",
  1136 => x"fefe4973",
  1137 => x"87e9f487",
  1138 => x"711e731e",
  1139 => x"4aa3c64b",
  1140 => x"c187dc02",
  1141 => x"e4c0028a",
  1142 => x"c1028a87",
  1143 => x"028a87e8",
  1144 => x"8a87cac1",
  1145 => x"87efc002",
  1146 => x"87d9028a",
  1147 => x"c287e9c1",
  1148 => x"df48e8ef",
  1149 => x"d549c178",
  1150 => x"e6c187ed",
  1151 => x"fc49c787",
  1152 => x"dec187f1",
  1153 => x"ecefc287",
  1154 => x"cbc102bf",
  1155 => x"88c14887",
  1156 => x"58f0efc2",
  1157 => x"c287c1c1",
  1158 => x"02bff0ef",
  1159 => x"c287f9c0",
  1160 => x"48bfecef",
  1161 => x"efc280c1",
  1162 => x"ebc058f0",
  1163 => x"ecefc287",
  1164 => x"89c649bf",
  1165 => x"59f0efc2",
  1166 => x"03a9b7c0",
  1167 => x"efc287da",
  1168 => x"78c048ec",
  1169 => x"efc287d2",
  1170 => x"cb02bff0",
  1171 => x"ecefc287",
  1172 => x"80c648bf",
  1173 => x"58f0efc2",
  1174 => x"cad449c0",
  1175 => x"c0497387",
  1176 => x"f287d4f9",
  1177 => x"5e0e87cb",
  1178 => x"710e5c5b",
  1179 => x"1e66cc4c",
  1180 => x"93cb4b74",
  1181 => x"83e0e1c1",
  1182 => x"6a4aa3c4",
  1183 => x"d1f9fe49",
  1184 => x"f1c3c187",
  1185 => x"49a3c87b",
  1186 => x"c95166d4",
  1187 => x"66d849a3",
  1188 => x"49a3ca51",
  1189 => x"265166dc",
  1190 => x"0e87d4f1",
  1191 => x"5d5c5b5e",
  1192 => x"86d0ff0e",
  1193 => x"c859a6d8",
  1194 => x"78c048a6",
  1195 => x"c4c180fc",
  1196 => x"80c87866",
  1197 => x"80c478c1",
  1198 => x"efc278c1",
  1199 => x"78c148f0",
  1200 => x"bfe8efc2",
  1201 => x"de486e7e",
  1202 => x"87cb05a8",
  1203 => x"7087d4f3",
  1204 => x"59a6cc49",
  1205 => x"6e87f8d0",
  1206 => x"05a8df48",
  1207 => x"c187eec1",
  1208 => x"c44966c0",
  1209 => x"c17e6981",
  1210 => x"6e48c4dd",
  1211 => x"4aa1d049",
  1212 => x"aa714120",
  1213 => x"c187f905",
  1214 => x"c14af1c3",
  1215 => x"7a0a66c0",
  1216 => x"66c0c10a",
  1217 => x"df81c949",
  1218 => x"66c0c151",
  1219 => x"c181ca49",
  1220 => x"c0c151d3",
  1221 => x"81cb4966",
  1222 => x"c44ba1c4",
  1223 => x"786b48a6",
  1224 => x"1e721e71",
  1225 => x"48d4ddc1",
  1226 => x"d04966cc",
  1227 => x"41204aa1",
  1228 => x"f905aa71",
  1229 => x"264a2687",
  1230 => x"c9797249",
  1231 => x"52df4aa1",
  1232 => x"d4c181ca",
  1233 => x"48a6c851",
  1234 => x"c2cf78c2",
  1235 => x"87ece587",
  1236 => x"e587cee6",
  1237 => x"4c7087db",
  1238 => x"02acfbc0",
  1239 => x"d487d0c1",
  1240 => x"c2c10566",
  1241 => x"1e1ec087",
  1242 => x"e3c11ec1",
  1243 => x"49c01ec3",
  1244 => x"c187f3fb",
  1245 => x"c44a66d0",
  1246 => x"c7496a82",
  1247 => x"c1517481",
  1248 => x"6a1ed81e",
  1249 => x"e581c849",
  1250 => x"86d887eb",
  1251 => x"4866c4c1",
  1252 => x"c701a8c0",
  1253 => x"48a6c887",
  1254 => x"87ce78c1",
  1255 => x"4866c4c1",
  1256 => x"a6c888c1",
  1257 => x"e487c358",
  1258 => x"a6cc87f7",
  1259 => x"7478c248",
  1260 => x"d6cd029c",
  1261 => x"4866c887",
  1262 => x"a866c8c1",
  1263 => x"87cbcd03",
  1264 => x"c048a6d8",
  1265 => x"87e9e378",
  1266 => x"d0c14c70",
  1267 => x"d6c205ac",
  1268 => x"7e66d887",
  1269 => x"7087cde6",
  1270 => x"59a6dc49",
  1271 => x"7087d2e3",
  1272 => x"acecc04c",
  1273 => x"87eac105",
  1274 => x"cb4966c8",
  1275 => x"66c0c191",
  1276 => x"4aa1c481",
  1277 => x"a1c84d6a",
  1278 => x"5266d84a",
  1279 => x"79f3c4c1",
  1280 => x"7087eee2",
  1281 => x"d8029c4c",
  1282 => x"acfbc087",
  1283 => x"7487d202",
  1284 => x"87dde255",
  1285 => x"029c4c70",
  1286 => x"fbc087c7",
  1287 => x"eeff05ac",
  1288 => x"55e0c087",
  1289 => x"c055c1c2",
  1290 => x"66d47d97",
  1291 => x"05a96e49",
  1292 => x"66c887db",
  1293 => x"a866c448",
  1294 => x"c887ca04",
  1295 => x"80c14866",
  1296 => x"c858a6cc",
  1297 => x"4866c487",
  1298 => x"a6c888c1",
  1299 => x"87e1e158",
  1300 => x"d0c14c70",
  1301 => x"87c805ac",
  1302 => x"c14866d0",
  1303 => x"58a6d480",
  1304 => x"02acd0c1",
  1305 => x"dc87eafd",
  1306 => x"66d448a6",
  1307 => x"4866d878",
  1308 => x"05a866dc",
  1309 => x"c087e6c9",
  1310 => x"c048a6e0",
  1311 => x"80c478f0",
  1312 => x"c47866cc",
  1313 => x"7e78c080",
  1314 => x"fbc04874",
  1315 => x"a6f0c088",
  1316 => x"02987058",
  1317 => x"4887e1c8",
  1318 => x"f0c088cb",
  1319 => x"987058a6",
  1320 => x"87e9c002",
  1321 => x"c088c948",
  1322 => x"7058a6f0",
  1323 => x"e9c30298",
  1324 => x"88c44887",
  1325 => x"58a6f0c0",
  1326 => x"d6029870",
  1327 => x"88c14887",
  1328 => x"58a6f0c0",
  1329 => x"c3029870",
  1330 => x"e5c787d0",
  1331 => x"a6e0c087",
  1332 => x"cc78c048",
  1333 => x"80c14866",
  1334 => x"ff58a6d0",
  1335 => x"7087d2df",
  1336 => x"acecc04c",
  1337 => x"c087d702",
  1338 => x"c00266e0",
  1339 => x"e4c087c7",
  1340 => x"c9c05ca6",
  1341 => x"c0487487",
  1342 => x"e8c088f0",
  1343 => x"ecc058a6",
  1344 => x"cdc002ac",
  1345 => x"e8deff87",
  1346 => x"c04c7087",
  1347 => x"ff05acec",
  1348 => x"e0c087f3",
  1349 => x"66d41e66",
  1350 => x"ecc01e49",
  1351 => x"e3c11e66",
  1352 => x"66d81ec3",
  1353 => x"87fef449",
  1354 => x"1eca1ec0",
  1355 => x"4966e0c0",
  1356 => x"d8c191cb",
  1357 => x"a6d88166",
  1358 => x"78a1c448",
  1359 => x"49bf66d8",
  1360 => x"87f1deff",
  1361 => x"b7c086d8",
  1362 => x"c8c106a8",
  1363 => x"de1ec187",
  1364 => x"bf66c81e",
  1365 => x"dcdeff49",
  1366 => x"7086c887",
  1367 => x"08c04849",
  1368 => x"a6e4c088",
  1369 => x"a8b7c058",
  1370 => x"87e9c006",
  1371 => x"4866e0c0",
  1372 => x"03a8b7dd",
  1373 => x"bf6e87df",
  1374 => x"66e0c049",
  1375 => x"51e0c081",
  1376 => x"81c14966",
  1377 => x"c281bf6e",
  1378 => x"e0c051c1",
  1379 => x"81c24966",
  1380 => x"c081bf6e",
  1381 => x"c47ec151",
  1382 => x"dfff87de",
  1383 => x"e4c087c6",
  1384 => x"deff58a6",
  1385 => x"e8c087fe",
  1386 => x"ecc058a6",
  1387 => x"cbc005a8",
  1388 => x"a6e4c087",
  1389 => x"66e0c048",
  1390 => x"87c4c078",
  1391 => x"87f1dbff",
  1392 => x"cb4966c8",
  1393 => x"66c0c191",
  1394 => x"70807148",
  1395 => x"c84a6e7e",
  1396 => x"ca496e82",
  1397 => x"66e0c081",
  1398 => x"66e4c051",
  1399 => x"c081c149",
  1400 => x"c18966e0",
  1401 => x"70307148",
  1402 => x"7189c149",
  1403 => x"f3c27a97",
  1404 => x"c049bfdd",
  1405 => x"972966e0",
  1406 => x"71484a6a",
  1407 => x"a6f0c098",
  1408 => x"c4496e58",
  1409 => x"dc4d6981",
  1410 => x"66d84866",
  1411 => x"c8c002a8",
  1412 => x"48a6d887",
  1413 => x"c5c078c0",
  1414 => x"48a6d887",
  1415 => x"66d878c1",
  1416 => x"1ee0c01e",
  1417 => x"dbff4975",
  1418 => x"86c887cb",
  1419 => x"b7c04c70",
  1420 => x"d4c106ac",
  1421 => x"c0857487",
  1422 => x"897449e0",
  1423 => x"ddc14b75",
  1424 => x"fe714ae4",
  1425 => x"c287fbe9",
  1426 => x"66e8c085",
  1427 => x"c080c148",
  1428 => x"c058a6ec",
  1429 => x"c14966ec",
  1430 => x"02a97081",
  1431 => x"d887c8c0",
  1432 => x"78c048a6",
  1433 => x"d887c5c0",
  1434 => x"78c148a6",
  1435 => x"c21e66d8",
  1436 => x"e0c049a4",
  1437 => x"70887148",
  1438 => x"49751e49",
  1439 => x"87f5d9ff",
  1440 => x"b7c086c8",
  1441 => x"c0ff01a8",
  1442 => x"66e8c087",
  1443 => x"87d1c002",
  1444 => x"81c9496e",
  1445 => x"5166e8c0",
  1446 => x"c6c1486e",
  1447 => x"ccc078c3",
  1448 => x"c9496e87",
  1449 => x"6e51c281",
  1450 => x"f7c6c148",
  1451 => x"c07ec178",
  1452 => x"d8ff87c6",
  1453 => x"4c7087eb",
  1454 => x"f5c0026e",
  1455 => x"4866c887",
  1456 => x"04a866c4",
  1457 => x"c887cbc0",
  1458 => x"80c14866",
  1459 => x"c058a6cc",
  1460 => x"66c487e0",
  1461 => x"c888c148",
  1462 => x"d5c058a6",
  1463 => x"acc6c187",
  1464 => x"87c8c005",
  1465 => x"c14866cc",
  1466 => x"58a6d080",
  1467 => x"87f1d7ff",
  1468 => x"66d04c70",
  1469 => x"d480c148",
  1470 => x"9c7458a6",
  1471 => x"87cbc002",
  1472 => x"c14866c8",
  1473 => x"04a866c8",
  1474 => x"ff87f5f2",
  1475 => x"c887c9d7",
  1476 => x"a8c74866",
  1477 => x"87e5c003",
  1478 => x"48f0efc2",
  1479 => x"66c878c0",
  1480 => x"c191cb49",
  1481 => x"c48166c0",
  1482 => x"4a6a4aa1",
  1483 => x"c87952c0",
  1484 => x"80c14866",
  1485 => x"c758a6cc",
  1486 => x"dbff04a8",
  1487 => x"8ed0ff87",
  1488 => x"87e9deff",
  1489 => x"64616f4c",
  1490 => x"74655320",
  1491 => x"676e6974",
  1492 => x"00812073",
  1493 => x"65766153",
  1494 => x"74655320",
  1495 => x"676e6974",
  1496 => x"00812073",
  1497 => x"1e00203a",
  1498 => x"4b711e73",
  1499 => x"87c6029b",
  1500 => x"48ecefc2",
  1501 => x"1ec778c0",
  1502 => x"bfecefc2",
  1503 => x"e1c11e49",
  1504 => x"efc21ee0",
  1505 => x"ec49bfe8",
  1506 => x"86cc87d1",
  1507 => x"bfe8efc2",
  1508 => x"87c7e749",
  1509 => x"c8029b73",
  1510 => x"e0e1c187",
  1511 => x"e8e5c049",
  1512 => x"ccddff87",
  1513 => x"f9c71e87",
  1514 => x"fe49c187",
  1515 => x"ecfe87f9",
  1516 => x"987087d9",
  1517 => x"fe87cd02",
  1518 => x"7087d6f5",
  1519 => x"87c40298",
  1520 => x"87c24ac1",
  1521 => x"9a724ac0",
  1522 => x"c087ce05",
  1523 => x"f6dfc11e",
  1524 => x"c3f1c049",
  1525 => x"fe86c487",
  1526 => x"c11ec087",
  1527 => x"c049c1e0",
  1528 => x"c087f5f0",
  1529 => x"cac2c11e",
  1530 => x"c0497087",
  1531 => x"c387e9f0",
  1532 => x"8ef887ef",
  1533 => x"44534f26",
  1534 => x"69616620",
  1535 => x"2e64656c",
  1536 => x"6f6f4200",
  1537 => x"676e6974",
  1538 => x"002e2e2e",
  1539 => x"d4e8c01e",
  1540 => x"f6f3c087",
  1541 => x"2687f687",
  1542 => x"efc21e4f",
  1543 => x"78c048ec",
  1544 => x"48e8efc2",
  1545 => x"fcfd78c0",
  1546 => x"c087e187",
  1547 => x"204f2648",
  1548 => x"20202020",
  1549 => x"20202020",
  1550 => x"20202020",
  1551 => x"74697845",
  1552 => x"20202020",
  1553 => x"20202020",
  1554 => x"20202020",
  1555 => x"20800081",
  1556 => x"20202020",
  1557 => x"20202020",
  1558 => x"42202020",
  1559 => x"006b6361",
  1560 => x"00001133",
  1561 => x"00002c01",
  1562 => x"33000000",
  1563 => x"1f000011",
  1564 => x"0000002c",
  1565 => x"11330000",
  1566 => x"2c3d0000",
  1567 => x"00000000",
  1568 => x"00113300",
  1569 => x"002c5b00",
  1570 => x"00000000",
  1571 => x"00001133",
  1572 => x"00002c79",
  1573 => x"33000000",
  1574 => x"97000011",
  1575 => x"0000002c",
  1576 => x"11330000",
  1577 => x"2cb50000",
  1578 => x"00000000",
  1579 => x"00113300",
  1580 => x"00000000",
  1581 => x"00000000",
  1582 => x"000011c8",
  1583 => x"00000000",
  1584 => x"4c000000",
  1585 => x"2064616f",
  1586 => x"1e002e2a",
  1587 => x"c048f0fe",
  1588 => x"7909cd78",
  1589 => x"1e4f2609",
  1590 => x"bff0fe1e",
  1591 => x"2626487e",
  1592 => x"f0fe1e4f",
  1593 => x"2678c148",
  1594 => x"f0fe1e4f",
  1595 => x"2678c048",
  1596 => x"4a711e4f",
  1597 => x"265252c0",
  1598 => x"5b5e0e4f",
  1599 => x"f40e5d5c",
  1600 => x"974d7186",
  1601 => x"a5c17e6d",
  1602 => x"486c974c",
  1603 => x"6e58a6c8",
  1604 => x"a866c448",
  1605 => x"ff87c505",
  1606 => x"87e6c048",
  1607 => x"c287caff",
  1608 => x"6c9749a5",
  1609 => x"4ba3714b",
  1610 => x"974b6b97",
  1611 => x"486e7e6c",
  1612 => x"a6c880c1",
  1613 => x"cc98c758",
  1614 => x"977058a6",
  1615 => x"87e1fe7c",
  1616 => x"8ef44873",
  1617 => x"4c264d26",
  1618 => x"4f264b26",
  1619 => x"5c5b5e0e",
  1620 => x"7186f40e",
  1621 => x"4a66d84c",
  1622 => x"c29affc3",
  1623 => x"6c974ba4",
  1624 => x"49a17349",
  1625 => x"6c975172",
  1626 => x"c1486e7e",
  1627 => x"58a6c880",
  1628 => x"a6cc98c7",
  1629 => x"f4547058",
  1630 => x"87caff8e",
  1631 => x"e8fd1e1e",
  1632 => x"4abfe087",
  1633 => x"c0e0c049",
  1634 => x"87cb0299",
  1635 => x"f3c21e72",
  1636 => x"f7fe49d3",
  1637 => x"fc86c487",
  1638 => x"7e7087fd",
  1639 => x"2687c2fd",
  1640 => x"c21e4f26",
  1641 => x"fd49d3f3",
  1642 => x"e5c187c7",
  1643 => x"dafc49fc",
  1644 => x"87d9c587",
  1645 => x"5e0e4f26",
  1646 => x"0e5d5c5b",
  1647 => x"bff2f3c2",
  1648 => x"cae8c14a",
  1649 => x"724c49bf",
  1650 => x"fc4d71bc",
  1651 => x"4bc087db",
  1652 => x"99d04974",
  1653 => x"7587d502",
  1654 => x"7199d049",
  1655 => x"c11ec01e",
  1656 => x"734adcee",
  1657 => x"c0491282",
  1658 => x"86c887e4",
  1659 => x"832d2cc1",
  1660 => x"ff04abc8",
  1661 => x"e8fb87da",
  1662 => x"cae8c187",
  1663 => x"f2f3c248",
  1664 => x"4d2678bf",
  1665 => x"4b264c26",
  1666 => x"00004f26",
  1667 => x"ff1e0000",
  1668 => x"e1c848d0",
  1669 => x"48d4ff78",
  1670 => x"66c478c5",
  1671 => x"c387c302",
  1672 => x"66c878e0",
  1673 => x"ff87c602",
  1674 => x"f0c348d4",
  1675 => x"48d4ff78",
  1676 => x"d0ff7871",
  1677 => x"78e1c848",
  1678 => x"2678e0c0",
  1679 => x"5b5e0e4f",
  1680 => x"4c710e5c",
  1681 => x"49d3f3c2",
  1682 => x"7087eefa",
  1683 => x"aab7c04a",
  1684 => x"87e3c204",
  1685 => x"05aae0c3",
  1686 => x"ecc187c9",
  1687 => x"78c148c0",
  1688 => x"c387d4c2",
  1689 => x"c905aaf0",
  1690 => x"fcebc187",
  1691 => x"c178c148",
  1692 => x"ecc187f5",
  1693 => x"c702bfc0",
  1694 => x"c24b7287",
  1695 => x"87c2b3c0",
  1696 => x"9c744b72",
  1697 => x"c187d105",
  1698 => x"1ebffceb",
  1699 => x"bfc0ecc1",
  1700 => x"fd49721e",
  1701 => x"86c887f8",
  1702 => x"bffcebc1",
  1703 => x"87e0c002",
  1704 => x"b7c44973",
  1705 => x"edc19129",
  1706 => x"4a7381dc",
  1707 => x"92c29acf",
  1708 => x"307248c1",
  1709 => x"baff4a70",
  1710 => x"98694872",
  1711 => x"87db7970",
  1712 => x"b7c44973",
  1713 => x"edc19129",
  1714 => x"4a7381dc",
  1715 => x"92c29acf",
  1716 => x"307248c3",
  1717 => x"69484a70",
  1718 => x"c17970b0",
  1719 => x"c048c0ec",
  1720 => x"fcebc178",
  1721 => x"c278c048",
  1722 => x"f849d3f3",
  1723 => x"4a7087cb",
  1724 => x"03aab7c0",
  1725 => x"c087ddfd",
  1726 => x"87c8fc48",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"494a711e",
  1730 => x"2687f2fc",
  1731 => x"4ac01e4f",
  1732 => x"91c44972",
  1733 => x"81dcedc1",
  1734 => x"82c179c0",
  1735 => x"04aab7d0",
  1736 => x"4f2687ee",
  1737 => x"5c5b5e0e",
  1738 => x"4d710e5d",
  1739 => x"7587faf6",
  1740 => x"2ab7c44a",
  1741 => x"dcedc192",
  1742 => x"cf4c7582",
  1743 => x"6a94c29c",
  1744 => x"2b744b49",
  1745 => x"48c29bc3",
  1746 => x"4c703074",
  1747 => x"4874bcff",
  1748 => x"7a709871",
  1749 => x"7387caf6",
  1750 => x"87e6fa48",
  1751 => x"00000000",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"00000000",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"25261e16",
  1768 => x"3e3d362e",
  1769 => x"48d0ff1e",
  1770 => x"7178e1c8",
  1771 => x"08d4ff48",
  1772 => x"1e4f2678",
  1773 => x"c848d0ff",
  1774 => x"487178e1",
  1775 => x"7808d4ff",
  1776 => x"ff4866c4",
  1777 => x"267808d4",
  1778 => x"4a711e4f",
  1779 => x"1e4966c4",
  1780 => x"deff4972",
  1781 => x"48d0ff87",
  1782 => x"2678e0c0",
  1783 => x"711e4f26",
  1784 => x"aab7c24a",
  1785 => x"8287c303",
  1786 => x"82ce87c2",
  1787 => x"721e66c4",
  1788 => x"87d5ff49",
  1789 => x"1e4f2626",
  1790 => x"c34ad4ff",
  1791 => x"d0ff7aff",
  1792 => x"78e1c848",
  1793 => x"f3c27ade",
  1794 => x"497abfdd",
  1795 => x"7028c848",
  1796 => x"d048717a",
  1797 => x"717a7028",
  1798 => x"7028d848",
  1799 => x"48d0ff7a",
  1800 => x"2678e0c0",
  1801 => x"5b5e0e4f",
  1802 => x"710e5d5c",
  1803 => x"ddf3c24c",
  1804 => x"744b4dbf",
  1805 => x"9b66d02b",
  1806 => x"66d483c1",
  1807 => x"87c204ab",
  1808 => x"4a744bc0",
  1809 => x"724966d0",
  1810 => x"75b9ff31",
  1811 => x"72487399",
  1812 => x"484a7030",
  1813 => x"f3c2b071",
  1814 => x"dafe58e1",
  1815 => x"264d2687",
  1816 => x"264b264c",
  1817 => x"d0ff1e4f",
  1818 => x"78c9c848",
  1819 => x"d4ff4871",
  1820 => x"4f267808",
  1821 => x"494a711e",
  1822 => x"d0ff87eb",
  1823 => x"2678c848",
  1824 => x"1e731e4f",
  1825 => x"f3c24b71",
  1826 => x"c302bfed",
  1827 => x"87ebc287",
  1828 => x"c848d0ff",
  1829 => x"497378c9",
  1830 => x"ffb1e0c0",
  1831 => x"787148d4",
  1832 => x"48e1f3c2",
  1833 => x"66c878c0",
  1834 => x"c387c502",
  1835 => x"87c249ff",
  1836 => x"f3c249c0",
  1837 => x"66cc59e9",
  1838 => x"c587c602",
  1839 => x"c44ad5d5",
  1840 => x"ffffcf87",
  1841 => x"edf3c24a",
  1842 => x"edf3c25a",
  1843 => x"c478c148",
  1844 => x"264d2687",
  1845 => x"264b264c",
  1846 => x"5b5e0e4f",
  1847 => x"710e5d5c",
  1848 => x"e9f3c24a",
  1849 => x"9a724cbf",
  1850 => x"4987cb02",
  1851 => x"f1c191c8",
  1852 => x"83714bf7",
  1853 => x"f5c187c4",
  1854 => x"4dc04bf7",
  1855 => x"99744913",
  1856 => x"bfe5f3c2",
  1857 => x"48d4ffb9",
  1858 => x"b7c17871",
  1859 => x"b7c8852c",
  1860 => x"87e804ad",
  1861 => x"bfe1f3c2",
  1862 => x"c280c848",
  1863 => x"fe58e5f3",
  1864 => x"731e87ef",
  1865 => x"134b711e",
  1866 => x"cb029a4a",
  1867 => x"fe497287",
  1868 => x"4a1387e7",
  1869 => x"87f5059a",
  1870 => x"1e87dafe",
  1871 => x"bfe1f3c2",
  1872 => x"e1f3c249",
  1873 => x"78a1c148",
  1874 => x"a9b7c0c4",
  1875 => x"ff87db03",
  1876 => x"f3c248d4",
  1877 => x"c278bfe5",
  1878 => x"49bfe1f3",
  1879 => x"48e1f3c2",
  1880 => x"c478a1c1",
  1881 => x"04a9b7c0",
  1882 => x"d0ff87e5",
  1883 => x"c278c848",
  1884 => x"c048edf3",
  1885 => x"004f2678",
  1886 => x"00000000",
  1887 => x"00000000",
  1888 => x"5f5f0000",
  1889 => x"00000000",
  1890 => x"03000303",
  1891 => x"14000003",
  1892 => x"7f147f7f",
  1893 => x"0000147f",
  1894 => x"6b6b2e24",
  1895 => x"4c00123a",
  1896 => x"6c18366a",
  1897 => x"30003256",
  1898 => x"77594f7e",
  1899 => x"0040683a",
  1900 => x"03070400",
  1901 => x"00000000",
  1902 => x"633e1c00",
  1903 => x"00000041",
  1904 => x"3e634100",
  1905 => x"0800001c",
  1906 => x"1c1c3e2a",
  1907 => x"00082a3e",
  1908 => x"3e3e0808",
  1909 => x"00000808",
  1910 => x"60e08000",
  1911 => x"00000000",
  1912 => x"08080808",
  1913 => x"00000808",
  1914 => x"60600000",
  1915 => x"40000000",
  1916 => x"0c183060",
  1917 => x"00010306",
  1918 => x"4d597f3e",
  1919 => x"00003e7f",
  1920 => x"7f7f0604",
  1921 => x"00000000",
  1922 => x"59716342",
  1923 => x"0000464f",
  1924 => x"49496322",
  1925 => x"1800367f",
  1926 => x"7f13161c",
  1927 => x"0000107f",
  1928 => x"45456727",
  1929 => x"0000397d",
  1930 => x"494b7e3c",
  1931 => x"00003079",
  1932 => x"79710101",
  1933 => x"0000070f",
  1934 => x"49497f36",
  1935 => x"0000367f",
  1936 => x"69494f06",
  1937 => x"00001e3f",
  1938 => x"66660000",
  1939 => x"00000000",
  1940 => x"66e68000",
  1941 => x"00000000",
  1942 => x"14140808",
  1943 => x"00002222",
  1944 => x"14141414",
  1945 => x"00001414",
  1946 => x"14142222",
  1947 => x"00000808",
  1948 => x"59510302",
  1949 => x"3e00060f",
  1950 => x"555d417f",
  1951 => x"00001e1f",
  1952 => x"09097f7e",
  1953 => x"00007e7f",
  1954 => x"49497f7f",
  1955 => x"0000367f",
  1956 => x"41633e1c",
  1957 => x"00004141",
  1958 => x"63417f7f",
  1959 => x"00001c3e",
  1960 => x"49497f7f",
  1961 => x"00004141",
  1962 => x"09097f7f",
  1963 => x"00000101",
  1964 => x"49417f3e",
  1965 => x"00007a7b",
  1966 => x"08087f7f",
  1967 => x"00007f7f",
  1968 => x"7f7f4100",
  1969 => x"00000041",
  1970 => x"40406020",
  1971 => x"7f003f7f",
  1972 => x"361c087f",
  1973 => x"00004163",
  1974 => x"40407f7f",
  1975 => x"7f004040",
  1976 => x"060c067f",
  1977 => x"7f007f7f",
  1978 => x"180c067f",
  1979 => x"00007f7f",
  1980 => x"41417f3e",
  1981 => x"00003e7f",
  1982 => x"09097f7f",
  1983 => x"3e00060f",
  1984 => x"7f61417f",
  1985 => x"0000407e",
  1986 => x"19097f7f",
  1987 => x"0000667f",
  1988 => x"594d6f26",
  1989 => x"0000327b",
  1990 => x"7f7f0101",
  1991 => x"00000101",
  1992 => x"40407f3f",
  1993 => x"00003f7f",
  1994 => x"70703f0f",
  1995 => x"7f000f3f",
  1996 => x"3018307f",
  1997 => x"41007f7f",
  1998 => x"1c1c3663",
  1999 => x"01416336",
  2000 => x"7c7c0603",
  2001 => x"61010306",
  2002 => x"474d5971",
  2003 => x"00004143",
  2004 => x"417f7f00",
  2005 => x"01000041",
  2006 => x"180c0603",
  2007 => x"00406030",
  2008 => x"7f414100",
  2009 => x"0800007f",
  2010 => x"0603060c",
  2011 => x"8000080c",
  2012 => x"80808080",
  2013 => x"00008080",
  2014 => x"07030000",
  2015 => x"00000004",
  2016 => x"54547420",
  2017 => x"0000787c",
  2018 => x"44447f7f",
  2019 => x"0000387c",
  2020 => x"44447c38",
  2021 => x"00000044",
  2022 => x"44447c38",
  2023 => x"00007f7f",
  2024 => x"54547c38",
  2025 => x"0000185c",
  2026 => x"057f7e04",
  2027 => x"00000005",
  2028 => x"a4a4bc18",
  2029 => x"00007cfc",
  2030 => x"04047f7f",
  2031 => x"0000787c",
  2032 => x"7d3d0000",
  2033 => x"00000040",
  2034 => x"fd808080",
  2035 => x"0000007d",
  2036 => x"38107f7f",
  2037 => x"0000446c",
  2038 => x"7f3f0000",
  2039 => x"7c000040",
  2040 => x"0c180c7c",
  2041 => x"0000787c",
  2042 => x"04047c7c",
  2043 => x"0000787c",
  2044 => x"44447c38",
  2045 => x"0000387c",
  2046 => x"2424fcfc",
  2047 => x"0000183c",
  2048 => x"24243c18",
  2049 => x"0000fcfc",
  2050 => x"04047c7c",
  2051 => x"0000080c",
  2052 => x"54545c48",
  2053 => x"00002074",
  2054 => x"447f3f04",
  2055 => x"00000044",
  2056 => x"40407c3c",
  2057 => x"00007c7c",
  2058 => x"60603c1c",
  2059 => x"3c001c3c",
  2060 => x"6030607c",
  2061 => x"44003c7c",
  2062 => x"3810386c",
  2063 => x"0000446c",
  2064 => x"60e0bc1c",
  2065 => x"00001c3c",
  2066 => x"5c746444",
  2067 => x"0000444c",
  2068 => x"773e0808",
  2069 => x"00004141",
  2070 => x"7f7f0000",
  2071 => x"00000000",
  2072 => x"3e774141",
  2073 => x"02000808",
  2074 => x"02030101",
  2075 => x"7f000102",
  2076 => x"7f7f7f7f",
  2077 => x"08007f7f",
  2078 => x"3e1c1c08",
  2079 => x"7f7f7f3e",
  2080 => x"1c3e3e7f",
  2081 => x"0008081c",
  2082 => x"7c7c1810",
  2083 => x"00001018",
  2084 => x"7c7c3010",
  2085 => x"10001030",
  2086 => x"78606030",
  2087 => x"4200061e",
  2088 => x"3c183c66",
  2089 => x"78004266",
  2090 => x"c6c26a38",
  2091 => x"6000386c",
  2092 => x"00600000",
  2093 => x"0e006000",
  2094 => x"5d5c5b5e",
  2095 => x"4c711e0e",
  2096 => x"bffef3c2",
  2097 => x"c04bc04d",
  2098 => x"02ab741e",
  2099 => x"a6c487c7",
  2100 => x"c578c048",
  2101 => x"48a6c487",
  2102 => x"66c478c1",
  2103 => x"ee49731e",
  2104 => x"86c887df",
  2105 => x"ef49e0c0",
  2106 => x"a5c487ef",
  2107 => x"f0496a4a",
  2108 => x"c6f187f0",
  2109 => x"c185cb87",
  2110 => x"abb7c883",
  2111 => x"87c7ff04",
  2112 => x"264d2626",
  2113 => x"264b264c",
  2114 => x"4a711e4f",
  2115 => x"5ac2f4c2",
  2116 => x"48c2f4c2",
  2117 => x"fe4978c7",
  2118 => x"4f2687dd",
  2119 => x"711e731e",
  2120 => x"aab7c04a",
  2121 => x"c287d303",
  2122 => x"05bfedd1",
  2123 => x"4bc187c4",
  2124 => x"4bc087c2",
  2125 => x"5bf1d1c2",
  2126 => x"d1c287c4",
  2127 => x"d1c25af1",
  2128 => x"c14abfed",
  2129 => x"a2c0c19a",
  2130 => x"87e8ec49",
  2131 => x"d1c248fc",
  2132 => x"fe78bfed",
  2133 => x"711e87ef",
  2134 => x"1e66c44a",
  2135 => x"fde94972",
  2136 => x"4f262687",
  2137 => x"edd1c21e",
  2138 => x"d7e649bf",
  2139 => x"f6f3c287",
  2140 => x"78bfe848",
  2141 => x"48f2f3c2",
  2142 => x"c278bfec",
  2143 => x"4abff6f3",
  2144 => x"99ffc349",
  2145 => x"722ab7c8",
  2146 => x"c2b07148",
  2147 => x"2658fef3",
  2148 => x"5b5e0e4f",
  2149 => x"710e5d5c",
  2150 => x"87c8ff4b",
  2151 => x"48f1f3c2",
  2152 => x"497350c0",
  2153 => x"7087fde5",
  2154 => x"9cc24c49",
  2155 => x"cb49eecb",
  2156 => x"497087c3",
  2157 => x"f1f3c24d",
  2158 => x"c105bf97",
  2159 => x"66d087e2",
  2160 => x"faf3c249",
  2161 => x"d60599bf",
  2162 => x"4966d487",
  2163 => x"bff2f3c2",
  2164 => x"87cb0599",
  2165 => x"cbe54973",
  2166 => x"02987087",
  2167 => x"c187c1c1",
  2168 => x"87c0fe4c",
  2169 => x"d8ca4975",
  2170 => x"02987087",
  2171 => x"f3c287c6",
  2172 => x"50c148f1",
  2173 => x"97f1f3c2",
  2174 => x"e3c005bf",
  2175 => x"faf3c287",
  2176 => x"66d049bf",
  2177 => x"d6ff0599",
  2178 => x"f2f3c287",
  2179 => x"66d449bf",
  2180 => x"caff0599",
  2181 => x"e4497387",
  2182 => x"987087ca",
  2183 => x"87fffe05",
  2184 => x"dcfb4874",
  2185 => x"5b5e0e87",
  2186 => x"f40e5d5c",
  2187 => x"4c4dc086",
  2188 => x"c47ebfec",
  2189 => x"f3c248a6",
  2190 => x"c178bffe",
  2191 => x"c71ec01e",
  2192 => x"87cdfd49",
  2193 => x"987086c8",
  2194 => x"ff87cd02",
  2195 => x"87ccfb49",
  2196 => x"e349dac1",
  2197 => x"4dc187ce",
  2198 => x"97f1f3c2",
  2199 => x"87c302bf",
  2200 => x"c287cad5",
  2201 => x"4bbff6f3",
  2202 => x"bfedd1c2",
  2203 => x"87e9c005",
  2204 => x"e249fdc3",
  2205 => x"fac387ee",
  2206 => x"87e8e249",
  2207 => x"ffc34973",
  2208 => x"c01e7199",
  2209 => x"87cefb49",
  2210 => x"b7c84973",
  2211 => x"c11e7129",
  2212 => x"87c2fb49",
  2213 => x"fac586c8",
  2214 => x"faf3c287",
  2215 => x"029b4bbf",
  2216 => x"d1c287dd",
  2217 => x"c749bfe9",
  2218 => x"987087d7",
  2219 => x"c087c405",
  2220 => x"c287d24b",
  2221 => x"fcc649e0",
  2222 => x"edd1c287",
  2223 => x"c287c658",
  2224 => x"c048e9d1",
  2225 => x"c2497378",
  2226 => x"87cd0599",
  2227 => x"e149ebc3",
  2228 => x"497087d2",
  2229 => x"c20299c2",
  2230 => x"734cfb87",
  2231 => x"0599c149",
  2232 => x"f4c387cd",
  2233 => x"87fce049",
  2234 => x"99c24970",
  2235 => x"fa87c202",
  2236 => x"c849734c",
  2237 => x"87cd0599",
  2238 => x"e049f5c3",
  2239 => x"497087e6",
  2240 => x"d40299c2",
  2241 => x"c2f4c287",
  2242 => x"87c902bf",
  2243 => x"c288c148",
  2244 => x"c258c6f4",
  2245 => x"c14cff87",
  2246 => x"c449734d",
  2247 => x"87ce0599",
  2248 => x"ff49f2c3",
  2249 => x"7087fddf",
  2250 => x"0299c249",
  2251 => x"f4c287db",
  2252 => x"487ebfc2",
  2253 => x"03a8b7c7",
  2254 => x"486e87cb",
  2255 => x"f4c280c1",
  2256 => x"c2c058c6",
  2257 => x"c14cfe87",
  2258 => x"49fdc34d",
  2259 => x"87d4dfff",
  2260 => x"99c24970",
  2261 => x"c287d502",
  2262 => x"02bfc2f4",
  2263 => x"c287c9c0",
  2264 => x"c048c2f4",
  2265 => x"87c2c078",
  2266 => x"4dc14cfd",
  2267 => x"ff49fac3",
  2268 => x"7087f1de",
  2269 => x"0299c249",
  2270 => x"f4c287d9",
  2271 => x"c748bfc2",
  2272 => x"c003a8b7",
  2273 => x"f4c287c9",
  2274 => x"78c748c2",
  2275 => x"fc87c2c0",
  2276 => x"c04dc14c",
  2277 => x"c003acb7",
  2278 => x"66c487d1",
  2279 => x"82d8c14a",
  2280 => x"c6c0026a",
  2281 => x"744b6a87",
  2282 => x"c00f7349",
  2283 => x"1ef0c31e",
  2284 => x"f749dac1",
  2285 => x"86c887db",
  2286 => x"c0029870",
  2287 => x"a6c887e2",
  2288 => x"c2f4c248",
  2289 => x"66c878bf",
  2290 => x"c491cb49",
  2291 => x"80714866",
  2292 => x"bf6e7e70",
  2293 => x"87c8c002",
  2294 => x"c84bbf6e",
  2295 => x"0f734966",
  2296 => x"c0029d75",
  2297 => x"f4c287c8",
  2298 => x"f349bfc2",
  2299 => x"d1c287c9",
  2300 => x"c002bff1",
  2301 => x"c24987dd",
  2302 => x"987087c7",
  2303 => x"87d3c002",
  2304 => x"bfc2f4c2",
  2305 => x"87eff249",
  2306 => x"cff449c0",
  2307 => x"f1d1c287",
  2308 => x"f478c048",
  2309 => x"87e9f38e",
  2310 => x"5c5b5e0e",
  2311 => x"711e0e5d",
  2312 => x"fef3c24c",
  2313 => x"cdc149bf",
  2314 => x"d1c14da1",
  2315 => x"747e6981",
  2316 => x"87cf029c",
  2317 => x"744ba5c4",
  2318 => x"fef3c27b",
  2319 => x"c8f349bf",
  2320 => x"747b6e87",
  2321 => x"87c4059c",
  2322 => x"87c24bc0",
  2323 => x"49734bc1",
  2324 => x"d487c9f3",
  2325 => x"87c70266",
  2326 => x"7087da49",
  2327 => x"c087c24a",
  2328 => x"f5d1c24a",
  2329 => x"d8f2265a",
  2330 => x"00000087",
  2331 => x"00000000",
  2332 => x"00000000",
  2333 => x"4a711e00",
  2334 => x"49bfc8ff",
  2335 => x"2648a172",
  2336 => x"c8ff1e4f",
  2337 => x"c0fe89bf",
  2338 => x"c0c0c0c0",
  2339 => x"87c401a9",
  2340 => x"87c24ac0",
  2341 => x"48724ac1",
  2342 => x"5e0e4f26",
  2343 => x"0e5d5c5b",
  2344 => x"d4ff4b71",
  2345 => x"4866d04c",
  2346 => x"49d678c0",
  2347 => x"87f4dbff",
  2348 => x"6c7cffc3",
  2349 => x"99ffc349",
  2350 => x"c3494d71",
  2351 => x"e0c199f0",
  2352 => x"87cb05a9",
  2353 => x"6c7cffc3",
  2354 => x"d098c348",
  2355 => x"c3780866",
  2356 => x"4a6c7cff",
  2357 => x"c331c849",
  2358 => x"4a6c7cff",
  2359 => x"4972b271",
  2360 => x"ffc331c8",
  2361 => x"714a6c7c",
  2362 => x"c84972b2",
  2363 => x"7cffc331",
  2364 => x"b2714a6c",
  2365 => x"c048d0ff",
  2366 => x"9b7378e0",
  2367 => x"7287c202",
  2368 => x"2648757b",
  2369 => x"264c264d",
  2370 => x"1e4f264b",
  2371 => x"86f81e73",
  2372 => x"a6c81e76",
  2373 => x"87c2fe49",
  2374 => x"4b7086c4",
  2375 => x"a8c4486e",
  2376 => x"87efc203",
  2377 => x"f0c34a73",
  2378 => x"aad0c19a",
  2379 => x"c187c702",
  2380 => x"c205aae0",
  2381 => x"9bc387dd",
  2382 => x"c487d802",
  2383 => x"31c94966",
  2384 => x"66c41e71",
  2385 => x"c292d44a",
  2386 => x"7249c6f4",
  2387 => x"eed1fe81",
  2388 => x"c286c487",
  2389 => x"f6c005ab",
  2390 => x"1e496e87",
  2391 => x"ff49e3c0",
  2392 => x"d887e6d9",
  2393 => x"fbd8ff49",
  2394 => x"1ec0c887",
  2395 => x"49f6e2c2",
  2396 => x"87fcedfd",
  2397 => x"c048d0ff",
  2398 => x"e2c278e0",
  2399 => x"66cc1ef6",
  2400 => x"c292d44a",
  2401 => x"7249c6f4",
  2402 => x"efcffe81",
  2403 => x"c186cc87",
  2404 => x"fec005ab",
  2405 => x"49f2c187",
  2406 => x"87f3eafd",
  2407 => x"1ef6e2c2",
  2408 => x"d44a66c4",
  2409 => x"c6f4c292",
  2410 => x"fe817249",
  2411 => x"c487cace",
  2412 => x"c01e4966",
  2413 => x"d8ff49e3",
  2414 => x"49d787cf",
  2415 => x"87e4d7ff",
  2416 => x"c21ec0c8",
  2417 => x"fd49f6e2",
  2418 => x"cc87d4ec",
  2419 => x"48d0ff86",
  2420 => x"f878e0c0",
  2421 => x"87effc8e",
  2422 => x"5c5b5e0e",
  2423 => x"711e0e5d",
  2424 => x"4cd4ff4d",
  2425 => x"487e66d4",
  2426 => x"06a8b7c4",
  2427 => x"48c087c5",
  2428 => x"7587e6c1",
  2429 => x"d7defe49",
  2430 => x"c41e7587",
  2431 => x"93d44b66",
  2432 => x"83c6f4c2",
  2433 => x"c9fe4973",
  2434 => x"83c887d3",
  2435 => x"d0ff4b6b",
  2436 => x"78e1c848",
  2437 => x"48737cdd",
  2438 => x"7098ffc3",
  2439 => x"c849737c",
  2440 => x"c3487129",
  2441 => x"7c7098ff",
  2442 => x"29d04973",
  2443 => x"ffc34871",
  2444 => x"737c7098",
  2445 => x"7028d848",
  2446 => x"7c7cc07c",
  2447 => x"7c7c7c7c",
  2448 => x"7c7c7c7c",
  2449 => x"d0ff7c7c",
  2450 => x"78e0c048",
  2451 => x"dc1e66c4",
  2452 => x"f4d5ff49",
  2453 => x"7386c887",
  2454 => x"e6fa2648",
  2455 => x"5b5e0e87",
  2456 => x"1e0e5d5c",
  2457 => x"d4ff7e71",
  2458 => x"c21e6e4b",
  2459 => x"fe49d6f5",
  2460 => x"c487eac7",
  2461 => x"9d4d7086",
  2462 => x"87c3c302",
  2463 => x"bfdef5c2",
  2464 => x"fe496e4c",
  2465 => x"ff87c9dc",
  2466 => x"c5c848d0",
  2467 => x"7bd6c178",
  2468 => x"7b154ac0",
  2469 => x"e0c082c1",
  2470 => x"f504aab7",
  2471 => x"48d0ff87",
  2472 => x"c5c878c4",
  2473 => x"7bd3c178",
  2474 => x"78c47bc1",
  2475 => x"c1029c74",
  2476 => x"e2c287fc",
  2477 => x"c0c87ef6",
  2478 => x"b7c08c4d",
  2479 => x"87c603ac",
  2480 => x"4da4c0c8",
  2481 => x"efc24cc0",
  2482 => x"49bf97e7",
  2483 => x"d20299d0",
  2484 => x"c21ec087",
  2485 => x"fe49d6f5",
  2486 => x"c487dec9",
  2487 => x"4a497086",
  2488 => x"c287efc0",
  2489 => x"c21ef6e2",
  2490 => x"fe49d6f5",
  2491 => x"c487cac9",
  2492 => x"4a497086",
  2493 => x"c848d0ff",
  2494 => x"d4c178c5",
  2495 => x"bf976e7b",
  2496 => x"c1486e7b",
  2497 => x"c17e7080",
  2498 => x"f0ff058d",
  2499 => x"48d0ff87",
  2500 => x"9a7278c4",
  2501 => x"c087c505",
  2502 => x"87e5c048",
  2503 => x"f5c21ec1",
  2504 => x"c6fe49d6",
  2505 => x"86c487f2",
  2506 => x"fe059c74",
  2507 => x"d0ff87c4",
  2508 => x"78c5c848",
  2509 => x"c07bd3c1",
  2510 => x"c178c47b",
  2511 => x"c087c248",
  2512 => x"4d262648",
  2513 => x"4b264c26",
  2514 => x"5e0e4f26",
  2515 => x"710e5c5b",
  2516 => x"0266cc4b",
  2517 => x"4c87e8c0",
  2518 => x"028cf0c0",
  2519 => x"7487e8c0",
  2520 => x"028ac14a",
  2521 => x"8a87e0c0",
  2522 => x"8a87dc02",
  2523 => x"c087d802",
  2524 => x"c0028ae0",
  2525 => x"8ac187e3",
  2526 => x"87e4c002",
  2527 => x"7387e8c0",
  2528 => x"87d9fb49",
  2529 => x"7487e2c0",
  2530 => x"f949c01e",
  2531 => x"1e7487ca",
  2532 => x"c3f94973",
  2533 => x"d086c887",
  2534 => x"c1497387",
  2535 => x"87c987e9",
  2536 => x"d5c24973",
  2537 => x"c087c287",
  2538 => x"87d8fe48",
  2539 => x"e1c21e00",
  2540 => x"c149bfef",
  2541 => x"f3e1c2b9",
  2542 => x"48d4ff59",
  2543 => x"ff78ffc3",
  2544 => x"e1c848d0",
  2545 => x"48d4ff78",
  2546 => x"31c478c1",
  2547 => x"d0ff7871",
  2548 => x"78e0c048",
  2549 => x"711e4f26",
  2550 => x"49a2c44a",
  2551 => x"48ddf3c2",
  2552 => x"4969786a",
  2553 => x"e1c2b9c1",
  2554 => x"c0ff59f3",
  2555 => x"c6d0ff87",
  2556 => x"2648c187",
  2557 => x"4a711e4f",
  2558 => x"c249a2c4",
  2559 => x"7abfddf3",
  2560 => x"bfefe1c2",
  2561 => x"1e4f2679",
  2562 => x"c21e4a71",
  2563 => x"fe49d6f5",
  2564 => x"c487cac1",
  2565 => x"02987086",
  2566 => x"e2c287dc",
  2567 => x"f5c21ef6",
  2568 => x"c4fe49d6",
  2569 => x"86c487d3",
  2570 => x"c9029870",
  2571 => x"f6e2c287",
  2572 => x"87e2fe49",
  2573 => x"48c087c2",
  2574 => x"711e4f26",
  2575 => x"f5c21e4a",
  2576 => x"c0fe49d6",
  2577 => x"86c487d7",
  2578 => x"de029870",
  2579 => x"f6e2c287",
  2580 => x"87e1fe49",
  2581 => x"1ef6e2c2",
  2582 => x"49d6f5c2",
  2583 => x"87dcc4fe",
  2584 => x"987086c4",
  2585 => x"c187c402",
  2586 => x"c087c248",
  2587 => x"004f2648",
  2588 => x"1e000000",
  2589 => x"bfc0e2c2",
  2590 => x"87e1f749",
  2591 => x"4f2648c0",
  2592 => x"00002884",
  2593 => x"54534d41",
  2594 => x"20444152",
  2595 => x"004d4f52",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
