library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fcc0c387",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49fcc0c3",
    18 => x"48d8e9c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"d8e9c287",
    25 => x"d4e9c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"efc187f7",
    29 => x"e9c287ee",
    30 => x"e9c24dd8",
    31 => x"ad744cd8",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87d0048b",
    67 => x"02114812",
    68 => x"c34c87ca",
    69 => x"749c98df",
    70 => x"87eb0288",
    71 => x"4b264a26",
    72 => x"4f264c26",
    73 => x"8148731e",
    74 => x"c502a973",
    75 => x"05531287",
    76 => x"4f2687f6",
    77 => x"721e731e",
    78 => x"e7c0029a",
    79 => x"c148c087",
    80 => x"06a9724b",
    81 => x"827287d1",
    82 => x"7387c906",
    83 => x"01a97283",
    84 => x"87c387f4",
    85 => x"723ab2c1",
    86 => x"738903a9",
    87 => x"2ac10780",
    88 => x"87f3052b",
    89 => x"4f264b26",
    90 => x"c41e751e",
    91 => x"a1b7714d",
    92 => x"c1b9ff04",
    93 => x"07bdc381",
    94 => x"04a2b772",
    95 => x"82c1baff",
    96 => x"fe07bdc1",
    97 => x"2dc187ee",
    98 => x"c1b8ff04",
    99 => x"042d0780",
   100 => x"81c1b9ff",
   101 => x"264d2607",
   102 => x"1e731e4f",
   103 => x"66c84a71",
   104 => x"8bc1494b",
   105 => x"cf029971",
   106 => x"ff481287",
   107 => x"737808d4",
   108 => x"718bc149",
   109 => x"87f10599",
   110 => x"4f264b26",
   111 => x"5c5b5e0e",
   112 => x"ff4a710e",
   113 => x"66cc4cd4",
   114 => x"8bc1494b",
   115 => x"ce029971",
   116 => x"7cffc387",
   117 => x"4973526c",
   118 => x"99718bc1",
   119 => x"2687f205",
   120 => x"264b264c",
   121 => x"1e731e4f",
   122 => x"c34bd4ff",
   123 => x"4a6b7bff",
   124 => x"6b7bffc3",
   125 => x"7232c849",
   126 => x"7bffc3b1",
   127 => x"31c84a6b",
   128 => x"ffc3b271",
   129 => x"c8496b7b",
   130 => x"71b17232",
   131 => x"264b2648",
   132 => x"5b5e0e4f",
   133 => x"710e5d5c",
   134 => x"4cd4ff4d",
   135 => x"ffc34875",
   136 => x"c27c7098",
   137 => x"05bfd8e9",
   138 => x"66d087c8",
   139 => x"d430c948",
   140 => x"66d058a6",
   141 => x"7129d849",
   142 => x"98ffc348",
   143 => x"66d07c70",
   144 => x"7129d049",
   145 => x"98ffc348",
   146 => x"66d07c70",
   147 => x"7129c849",
   148 => x"98ffc348",
   149 => x"66d07c70",
   150 => x"98ffc348",
   151 => x"49757c70",
   152 => x"487129d0",
   153 => x"7098ffc3",
   154 => x"c94b6c7c",
   155 => x"c34afff0",
   156 => x"cf05abff",
   157 => x"7c714987",
   158 => x"8ac14b6c",
   159 => x"7187c502",
   160 => x"87f202ab",
   161 => x"4d264873",
   162 => x"4b264c26",
   163 => x"c01e4f26",
   164 => x"48d4ff49",
   165 => x"c178ffc3",
   166 => x"b7c8c381",
   167 => x"87f104a9",
   168 => x"5e0e4f26",
   169 => x"0e5d5c5b",
   170 => x"c1f0ffc0",
   171 => x"c0c14df7",
   172 => x"c0c0c0c0",
   173 => x"87d6ff4b",
   174 => x"4cdff8c4",
   175 => x"49751ec0",
   176 => x"c487cefd",
   177 => x"05a8c186",
   178 => x"ff87e5c0",
   179 => x"ffc348d4",
   180 => x"c01e7378",
   181 => x"e9c1f0e1",
   182 => x"87f5fc49",
   183 => x"987086c4",
   184 => x"ff87ca05",
   185 => x"ffc348d4",
   186 => x"cb48c178",
   187 => x"87defe87",
   188 => x"ff058cc1",
   189 => x"48c087c6",
   190 => x"4c264d26",
   191 => x"4f264b26",
   192 => x"5c5b5e0e",
   193 => x"f0ffc00e",
   194 => x"ff4cc1c1",
   195 => x"ffc348d4",
   196 => x"49c4cd78",
   197 => x"d387d0f6",
   198 => x"741ec04b",
   199 => x"87f1fb49",
   200 => x"987086c4",
   201 => x"ff87ca05",
   202 => x"ffc348d4",
   203 => x"cb48c178",
   204 => x"87dafd87",
   205 => x"ff058bc1",
   206 => x"48c087df",
   207 => x"4b264c26",
   208 => x"00004f26",
   209 => x"00444d43",
   210 => x"5c5b5e0e",
   211 => x"ffc30e5d",
   212 => x"4bd4ff4d",
   213 => x"c687f7fc",
   214 => x"e1c01eea",
   215 => x"49c8c1f0",
   216 => x"c487eefa",
   217 => x"02a8c186",
   218 => x"d3fe87c8",
   219 => x"c148c087",
   220 => x"f0f987e8",
   221 => x"cf497087",
   222 => x"c699ffff",
   223 => x"c802a9ea",
   224 => x"87fcfd87",
   225 => x"d1c148c0",
   226 => x"c07b7587",
   227 => x"d1fc4cf1",
   228 => x"02987087",
   229 => x"c087ecc0",
   230 => x"f0ffc01e",
   231 => x"f949fac1",
   232 => x"86c487ef",
   233 => x"da059870",
   234 => x"6b7b7587",
   235 => x"757b7549",
   236 => x"757b757b",
   237 => x"99c0c17b",
   238 => x"c187c402",
   239 => x"c087db48",
   240 => x"c287d748",
   241 => x"87ca05ac",
   242 => x"f349e4cf",
   243 => x"48c087d9",
   244 => x"8cc187c8",
   245 => x"87f6fe05",
   246 => x"4d2648c0",
   247 => x"4b264c26",
   248 => x"00004f26",
   249 => x"43484453",
   250 => x"69616620",
   251 => x"000a216c",
   252 => x"5c5b5e0e",
   253 => x"d0ff0e5d",
   254 => x"d0e5c04d",
   255 => x"c24cc0c1",
   256 => x"c148d8e9",
   257 => x"49fcd178",
   258 => x"c787dcf2",
   259 => x"f97dc24b",
   260 => x"7dc387fc",
   261 => x"49741ec0",
   262 => x"c487f6f7",
   263 => x"05a8c186",
   264 => x"c24b87c1",
   265 => x"87cb05ab",
   266 => x"f149f4d1",
   267 => x"48c087f9",
   268 => x"c187f6c0",
   269 => x"d4ff058b",
   270 => x"87ccfc87",
   271 => x"58dce9c2",
   272 => x"cd059870",
   273 => x"c01ec187",
   274 => x"d0c1f0ff",
   275 => x"87c1f749",
   276 => x"d4ff86c4",
   277 => x"78ffc348",
   278 => x"c287ccc5",
   279 => x"c258e0e9",
   280 => x"48d4ff7d",
   281 => x"c178ffc3",
   282 => x"264d2648",
   283 => x"264b264c",
   284 => x"0000004f",
   285 => x"52524549",
   286 => x"00000000",
   287 => x"00495053",
   288 => x"5c5b5e0e",
   289 => x"4d710e5d",
   290 => x"ff4cffc3",
   291 => x"7b744bd4",
   292 => x"c448d0ff",
   293 => x"7b7478c3",
   294 => x"ffc01e75",
   295 => x"49d8c1f0",
   296 => x"c487eef5",
   297 => x"02987086",
   298 => x"ecd387cb",
   299 => x"87f7ef49",
   300 => x"eec048c1",
   301 => x"c37b7487",
   302 => x"c0c87bfe",
   303 => x"4966d41e",
   304 => x"c487d6f3",
   305 => x"747b7486",
   306 => x"d87b747b",
   307 => x"744ae0da",
   308 => x"c5056b7b",
   309 => x"058ac187",
   310 => x"7b7487f5",
   311 => x"c248d0ff",
   312 => x"2648c078",
   313 => x"264c264d",
   314 => x"004f264b",
   315 => x"74697257",
   316 => x"61662065",
   317 => x"64656c69",
   318 => x"5e0e000a",
   319 => x"0e5d5c5b",
   320 => x"4b7186fc",
   321 => x"c04cd4ff",
   322 => x"cdeec57e",
   323 => x"ffc34adf",
   324 => x"c3486c7c",
   325 => x"c005a8fe",
   326 => x"4d7487f8",
   327 => x"cc029b73",
   328 => x"1e66d487",
   329 => x"d3f24973",
   330 => x"d486c487",
   331 => x"48d0ff87",
   332 => x"d478d1c4",
   333 => x"ffc34a66",
   334 => x"058ac17d",
   335 => x"a6d887f8",
   336 => x"7cffc35a",
   337 => x"059b737c",
   338 => x"d0ff87c5",
   339 => x"c178d048",
   340 => x"8ac17e4a",
   341 => x"87f6fe05",
   342 => x"8efc486e",
   343 => x"4c264d26",
   344 => x"4f264b26",
   345 => x"711e731e",
   346 => x"ff4bc04a",
   347 => x"ffc348d4",
   348 => x"48d0ff78",
   349 => x"ff78c3c4",
   350 => x"ffc348d4",
   351 => x"c01e7278",
   352 => x"d1c1f0ff",
   353 => x"87c9f249",
   354 => x"987086c4",
   355 => x"c887d205",
   356 => x"66cc1ec0",
   357 => x"87e2fd49",
   358 => x"4b7086c4",
   359 => x"c248d0ff",
   360 => x"26487378",
   361 => x"0e4f264b",
   362 => x"5d5c5b5e",
   363 => x"c01ec00e",
   364 => x"c9c1f0ff",
   365 => x"87d9f149",
   366 => x"e9c21ed2",
   367 => x"f9fc49e0",
   368 => x"c086c887",
   369 => x"d284c14c",
   370 => x"f804acb7",
   371 => x"e0e9c287",
   372 => x"c349bf97",
   373 => x"c0c199c0",
   374 => x"e7c005a9",
   375 => x"e7e9c287",
   376 => x"d049bf97",
   377 => x"e8e9c231",
   378 => x"c84abf97",
   379 => x"c2b17232",
   380 => x"bf97e9e9",
   381 => x"4c71b14a",
   382 => x"ffffffcf",
   383 => x"ca84c19c",
   384 => x"87e7c134",
   385 => x"97e9e9c2",
   386 => x"31c149bf",
   387 => x"e9c299c6",
   388 => x"4abf97ea",
   389 => x"722ab7c7",
   390 => x"e5e9c2b1",
   391 => x"4d4abf97",
   392 => x"e9c29dcf",
   393 => x"4abf97e6",
   394 => x"32ca9ac3",
   395 => x"97e7e9c2",
   396 => x"33c24bbf",
   397 => x"e9c2b273",
   398 => x"4bbf97e8",
   399 => x"c69bc0c3",
   400 => x"b2732bb7",
   401 => x"48c181c2",
   402 => x"49703071",
   403 => x"307548c1",
   404 => x"4c724d70",
   405 => x"947184c1",
   406 => x"adb7c0c8",
   407 => x"c187cc06",
   408 => x"c82db734",
   409 => x"01adb7c0",
   410 => x"7487f4ff",
   411 => x"264d2648",
   412 => x"264b264c",
   413 => x"5b5e0e4f",
   414 => x"f80e5d5c",
   415 => x"c8f2c286",
   416 => x"c278c048",
   417 => x"c01ec0ea",
   418 => x"87d8fb49",
   419 => x"987086c4",
   420 => x"c087c505",
   421 => x"87c0c948",
   422 => x"7ec14dc0",
   423 => x"bfc0ffc0",
   424 => x"f6eac249",
   425 => x"4bc8714a",
   426 => x"7087fbe8",
   427 => x"87c20598",
   428 => x"fec07ec0",
   429 => x"c249bffc",
   430 => x"714ad2eb",
   431 => x"e5e84bc8",
   432 => x"05987087",
   433 => x"7ec087c2",
   434 => x"fdc0026e",
   435 => x"c6f1c287",
   436 => x"f1c24dbf",
   437 => x"7ebf9ffe",
   438 => x"ead6c548",
   439 => x"87c705a8",
   440 => x"bfc6f1c2",
   441 => x"6e87ce4d",
   442 => x"d5e9ca48",
   443 => x"87c502a8",
   444 => x"e3c748c0",
   445 => x"c0eac287",
   446 => x"f949751e",
   447 => x"86c487e6",
   448 => x"c5059870",
   449 => x"c748c087",
   450 => x"fec087ce",
   451 => x"c249bffc",
   452 => x"714ad2eb",
   453 => x"cde74bc8",
   454 => x"05987087",
   455 => x"f2c287c8",
   456 => x"78c148c8",
   457 => x"ffc087da",
   458 => x"c249bfc0",
   459 => x"714af6ea",
   460 => x"f1e64bc8",
   461 => x"02987087",
   462 => x"c087c5c0",
   463 => x"87d8c648",
   464 => x"97fef1c2",
   465 => x"d5c149bf",
   466 => x"cdc005a9",
   467 => x"fff1c287",
   468 => x"c249bf97",
   469 => x"c002a9ea",
   470 => x"48c087c5",
   471 => x"c287f9c5",
   472 => x"bf97c0ea",
   473 => x"e9c3487e",
   474 => x"cec002a8",
   475 => x"c3486e87",
   476 => x"c002a8eb",
   477 => x"48c087c5",
   478 => x"c287ddc5",
   479 => x"bf97cbea",
   480 => x"c0059949",
   481 => x"eac287cc",
   482 => x"49bf97cc",
   483 => x"c002a9c2",
   484 => x"48c087c5",
   485 => x"c287c1c5",
   486 => x"bf97cdea",
   487 => x"c4f2c248",
   488 => x"484c7058",
   489 => x"f2c288c1",
   490 => x"eac258c8",
   491 => x"49bf97ce",
   492 => x"eac28175",
   493 => x"4abf97cf",
   494 => x"a17232c8",
   495 => x"d8f6c27e",
   496 => x"c2786e48",
   497 => x"bf97d0ea",
   498 => x"58a6c848",
   499 => x"bfc8f2c2",
   500 => x"87cfc202",
   501 => x"bffcfec0",
   502 => x"d2ebc249",
   503 => x"4bc8714a",
   504 => x"7087c3e4",
   505 => x"c5c00298",
   506 => x"c348c087",
   507 => x"f2c287ea",
   508 => x"c24cbfc0",
   509 => x"c25cecf6",
   510 => x"bf97e5ea",
   511 => x"c231c849",
   512 => x"bf97e4ea",
   513 => x"c249a14a",
   514 => x"bf97e6ea",
   515 => x"7232d04a",
   516 => x"eac249a1",
   517 => x"4abf97e7",
   518 => x"a17232d8",
   519 => x"9166c449",
   520 => x"bfd8f6c2",
   521 => x"e0f6c281",
   522 => x"edeac259",
   523 => x"c84abf97",
   524 => x"eceac232",
   525 => x"a24bbf97",
   526 => x"eeeac24a",
   527 => x"d04bbf97",
   528 => x"4aa27333",
   529 => x"97efeac2",
   530 => x"9bcf4bbf",
   531 => x"a27333d8",
   532 => x"e4f6c24a",
   533 => x"748ac25a",
   534 => x"e4f6c292",
   535 => x"78a17248",
   536 => x"c287c1c1",
   537 => x"bf97d2ea",
   538 => x"c231c849",
   539 => x"bf97d1ea",
   540 => x"c549a14a",
   541 => x"81ffc731",
   542 => x"f6c229c9",
   543 => x"eac259ec",
   544 => x"4abf97d7",
   545 => x"eac232c8",
   546 => x"4bbf97d6",
   547 => x"66c44aa2",
   548 => x"c2826e92",
   549 => x"c25ae8f6",
   550 => x"c048e0f6",
   551 => x"dcf6c278",
   552 => x"78a17248",
   553 => x"48ecf6c2",
   554 => x"bfe0f6c2",
   555 => x"f0f6c278",
   556 => x"e4f6c248",
   557 => x"f2c278bf",
   558 => x"c002bfc8",
   559 => x"487487c9",
   560 => x"7e7030c4",
   561 => x"c287c9c0",
   562 => x"48bfe8f6",
   563 => x"7e7030c4",
   564 => x"48ccf2c2",
   565 => x"48c1786e",
   566 => x"4d268ef8",
   567 => x"4b264c26",
   568 => x"5e0e4f26",
   569 => x"0e5d5c5b",
   570 => x"f2c24a71",
   571 => x"cb02bfc8",
   572 => x"c74b7287",
   573 => x"c14d722b",
   574 => x"87c99dff",
   575 => x"2bc84b72",
   576 => x"ffc34d72",
   577 => x"d8f6c29d",
   578 => x"fec083bf",
   579 => x"02abbff8",
   580 => x"fec087d9",
   581 => x"eac25bfc",
   582 => x"49731ec0",
   583 => x"c487c5f1",
   584 => x"05987086",
   585 => x"48c087c5",
   586 => x"c287e6c0",
   587 => x"02bfc8f2",
   588 => x"497587d2",
   589 => x"eac291c4",
   590 => x"4c6981c0",
   591 => x"ffffffcf",
   592 => x"87cb9cff",
   593 => x"91c24975",
   594 => x"81c0eac2",
   595 => x"744c699f",
   596 => x"264d2648",
   597 => x"264b264c",
   598 => x"5b5e0e4f",
   599 => x"f00e5d5c",
   600 => x"59a6cc86",
   601 => x"c50566c8",
   602 => x"c448c087",
   603 => x"66c887c4",
   604 => x"7080c848",
   605 => x"78c0487e",
   606 => x"0266e0c0",
   607 => x"e0c087c8",
   608 => x"05bf9766",
   609 => x"48c087c5",
   610 => x"c087e7c3",
   611 => x"4949c11e",
   612 => x"c487ead0",
   613 => x"9c4c7086",
   614 => x"87fec002",
   615 => x"4ad0f2c2",
   616 => x"4966e0c0",
   617 => x"87e3dcff",
   618 => x"c0029870",
   619 => x"4a7487ec",
   620 => x"4966e0c0",
   621 => x"ddff4bcb",
   622 => x"987087c6",
   623 => x"c087db02",
   624 => x"029c741e",
   625 => x"4dc087c4",
   626 => x"4dc187c2",
   627 => x"eccf4975",
   628 => x"7086c487",
   629 => x"ff059c4c",
   630 => x"9c7487c2",
   631 => x"87d0c202",
   632 => x"6e49a4dc",
   633 => x"da786948",
   634 => x"66c849a4",
   635 => x"c880c448",
   636 => x"699f58a6",
   637 => x"0866c448",
   638 => x"c8f2c278",
   639 => x"87d202bf",
   640 => x"9f49a4d4",
   641 => x"ffc04969",
   642 => x"487199ff",
   643 => x"58a630d0",
   644 => x"a6cc87c5",
   645 => x"cc78c048",
   646 => x"66c44866",
   647 => x"66c480bf",
   648 => x"66c87808",
   649 => x"c878c048",
   650 => x"81cc4966",
   651 => x"79bf66c4",
   652 => x"d04966c8",
   653 => x"4d79c081",
   654 => x"c84c66c4",
   655 => x"82d44a66",
   656 => x"91c84975",
   657 => x"c049a172",
   658 => x"c1796c41",
   659 => x"adb7c685",
   660 => x"87e7ff04",
   661 => x"c94abf6e",
   662 => x"c049722a",
   663 => x"dbff4af0",
   664 => x"4a7087d2",
   665 => x"c14966c8",
   666 => x"797281c4",
   667 => x"87c248c1",
   668 => x"8ef048c0",
   669 => x"4c264d26",
   670 => x"4f264b26",
   671 => x"5c5b5e0e",
   672 => x"4c710e5d",
   673 => x"744d66d0",
   674 => x"c2c1029c",
   675 => x"49a4c887",
   676 => x"fac00269",
   677 => x"85496c87",
   678 => x"f2c2b975",
   679 => x"ff4abfc4",
   680 => x"719972ba",
   681 => x"e4c00299",
   682 => x"4ba4c487",
   683 => x"f1f8496b",
   684 => x"c27b7087",
   685 => x"49bfc0f2",
   686 => x"7c71816c",
   687 => x"f2c2b975",
   688 => x"ff4abfc4",
   689 => x"719972ba",
   690 => x"dcff0599",
   691 => x"267c7587",
   692 => x"264c264d",
   693 => x"1e4f264b",
   694 => x"4b711e73",
   695 => x"87c7029b",
   696 => x"6949a3c8",
   697 => x"c087c505",
   698 => x"87f6c048",
   699 => x"bfdcf6c2",
   700 => x"4aa3c449",
   701 => x"8ac24a6a",
   702 => x"bfc0f2c2",
   703 => x"49a17292",
   704 => x"bfc4f2c2",
   705 => x"729a6b4a",
   706 => x"fec049a1",
   707 => x"66c859fc",
   708 => x"cfe9711e",
   709 => x"7086c487",
   710 => x"87c40598",
   711 => x"87c248c0",
   712 => x"4b2648c1",
   713 => x"731e4f26",
   714 => x"9b4b711e",
   715 => x"c887c702",
   716 => x"056949a3",
   717 => x"48c087c5",
   718 => x"c287f6c0",
   719 => x"49bfdcf6",
   720 => x"6a4aa3c4",
   721 => x"c28ac24a",
   722 => x"92bfc0f2",
   723 => x"c249a172",
   724 => x"4abfc4f2",
   725 => x"a1729a6b",
   726 => x"fcfec049",
   727 => x"1e66c859",
   728 => x"87dce471",
   729 => x"987086c4",
   730 => x"c087c405",
   731 => x"c187c248",
   732 => x"264b2648",
   733 => x"5b5e0e4f",
   734 => x"f80e5d5c",
   735 => x"c47e7186",
   736 => x"78ff48a6",
   737 => x"ffffffc1",
   738 => x"c04dffff",
   739 => x"d44a6e4b",
   740 => x"c8497382",
   741 => x"49a17291",
   742 => x"694c66d8",
   743 => x"acb7c08c",
   744 => x"7587cb04",
   745 => x"c503acb7",
   746 => x"5ba6c887",
   747 => x"83c14d74",
   748 => x"04abb7c6",
   749 => x"c487d6ff",
   750 => x"8ef84866",
   751 => x"4c264d26",
   752 => x"4f264b26",
   753 => x"5c5b5e0e",
   754 => x"86f00e5d",
   755 => x"a6c47e71",
   756 => x"ffffc148",
   757 => x"78ffffff",
   758 => x"78ff80c4",
   759 => x"4cc04dc0",
   760 => x"83d44b6e",
   761 => x"92c84a74",
   762 => x"754aa273",
   763 => x"7391c849",
   764 => x"486a49a1",
   765 => x"49708869",
   766 => x"7459a6d0",
   767 => x"87d202ad",
   768 => x"c44866cc",
   769 => x"c903a866",
   770 => x"5ca6cc87",
   771 => x"cc48a6c4",
   772 => x"84c17866",
   773 => x"04acb7c6",
   774 => x"c187c5ff",
   775 => x"adb7c685",
   776 => x"87fafe04",
   777 => x"f04866c8",
   778 => x"264d268e",
   779 => x"264b264c",
   780 => x"5b5e0e4f",
   781 => x"ec0e5d5c",
   782 => x"c04b7186",
   783 => x"c94866e4",
   784 => x"58a6c828",
   785 => x"bfc4f2c2",
   786 => x"72baff4a",
   787 => x"9866c448",
   788 => x"7358a6cc",
   789 => x"c1c3029b",
   790 => x"49a3c887",
   791 => x"f9c20269",
   792 => x"6b487287",
   793 => x"58a6d498",
   794 => x"6c4ca3c4",
   795 => x"4866c87e",
   796 => x"05a866d0",
   797 => x"66c487c6",
   798 => x"87ccc27b",
   799 => x"731e66c8",
   800 => x"87f1fb49",
   801 => x"4d7086c4",
   802 => x"04adb7c0",
   803 => x"a3d487d0",
   804 => x"c849754a",
   805 => x"49a17291",
   806 => x"7c697b21",
   807 => x"7bc087c7",
   808 => x"6949a3cc",
   809 => x"4866c47c",
   810 => x"a6c8886b",
   811 => x"1e66d058",
   812 => x"c0fb4973",
   813 => x"7086c487",
   814 => x"a3c4c14d",
   815 => x"48a6c849",
   816 => x"66d07869",
   817 => x"a866c848",
   818 => x"87f2c006",
   819 => x"04adb7c0",
   820 => x"cc87ebc0",
   821 => x"a3d448a6",
   822 => x"c8497578",
   823 => x"8166cc91",
   824 => x"694866d0",
   825 => x"c8497088",
   826 => x"d106a966",
   827 => x"fb497387",
   828 => x"497087d2",
   829 => x"66cc91c8",
   830 => x"4166d081",
   831 => x"66c4796e",
   832 => x"f549731e",
   833 => x"86c487f6",
   834 => x"1ec0eac2",
   835 => x"c6f74973",
   836 => x"d086c487",
   837 => x"e4c049a3",
   838 => x"8eec7966",
   839 => x"4c264d26",
   840 => x"4f264b26",
   841 => x"711e731e",
   842 => x"c0029b4b",
   843 => x"f6c287e4",
   844 => x"4a735bf0",
   845 => x"f2c28ac2",
   846 => x"9249bfc0",
   847 => x"bfdcf6c2",
   848 => x"c2807248",
   849 => x"7158f4f6",
   850 => x"c230c448",
   851 => x"c058d0f2",
   852 => x"f6c287ed",
   853 => x"f6c248ec",
   854 => x"c278bfe0",
   855 => x"c248f0f6",
   856 => x"78bfe4f6",
   857 => x"bfc8f2c2",
   858 => x"c287c902",
   859 => x"49bfc0f2",
   860 => x"87c731c4",
   861 => x"bfe8f6c2",
   862 => x"c231c449",
   863 => x"2659d0f2",
   864 => x"0e4f264b",
   865 => x"0e5c5b5e",
   866 => x"4bc04a71",
   867 => x"c0029a72",
   868 => x"a2da87e0",
   869 => x"4b699f49",
   870 => x"bfc8f2c2",
   871 => x"d487cf02",
   872 => x"699f49a2",
   873 => x"ffc04c49",
   874 => x"34d09cff",
   875 => x"4cc087c2",
   876 => x"4973b374",
   877 => x"2687edfd",
   878 => x"264b264c",
   879 => x"5b5e0e4f",
   880 => x"f00e5d5c",
   881 => x"59a6c886",
   882 => x"ffffffcf",
   883 => x"7ec04cf8",
   884 => x"d80266c4",
   885 => x"fce9c287",
   886 => x"c278c048",
   887 => x"c248f4e9",
   888 => x"78bff0f6",
   889 => x"48f8e9c2",
   890 => x"bfecf6c2",
   891 => x"ddf2c278",
   892 => x"c250c048",
   893 => x"49bfccf2",
   894 => x"bffce9c2",
   895 => x"03aa714a",
   896 => x"7287ccc4",
   897 => x"0599cf49",
   898 => x"c087eac0",
   899 => x"c248f8fe",
   900 => x"78bff4e9",
   901 => x"1ec0eac2",
   902 => x"bff4e9c2",
   903 => x"f4e9c249",
   904 => x"78a1c148",
   905 => x"fbdcff71",
   906 => x"c086c487",
   907 => x"c248f4fe",
   908 => x"cc78c0ea",
   909 => x"f4fec087",
   910 => x"e0c048bf",
   911 => x"f8fec080",
   912 => x"fce9c258",
   913 => x"80c148bf",
   914 => x"58c0eac2",
   915 => x"000fb427",
   916 => x"bf97bf00",
   917 => x"c2029d4d",
   918 => x"e5c387e5",
   919 => x"dec202ad",
   920 => x"f4fec087",
   921 => x"a3cb4bbf",
   922 => x"cf4c1149",
   923 => x"d2c105ac",
   924 => x"df497587",
   925 => x"cd89c199",
   926 => x"d0f2c291",
   927 => x"4aa3c181",
   928 => x"a3c35112",
   929 => x"c551124a",
   930 => x"51124aa3",
   931 => x"124aa3c7",
   932 => x"4aa3c951",
   933 => x"a3ce5112",
   934 => x"d051124a",
   935 => x"51124aa3",
   936 => x"124aa3d2",
   937 => x"4aa3d451",
   938 => x"a3d65112",
   939 => x"d851124a",
   940 => x"51124aa3",
   941 => x"124aa3dc",
   942 => x"4aa3de51",
   943 => x"7ec15112",
   944 => x"7487fcc0",
   945 => x"0599c849",
   946 => x"7487edc0",
   947 => x"0599d049",
   948 => x"e0c087d3",
   949 => x"ccc00266",
   950 => x"c0497387",
   951 => x"700f66e0",
   952 => x"d3c00298",
   953 => x"c0056e87",
   954 => x"f2c287c6",
   955 => x"50c048d0",
   956 => x"bff4fec0",
   957 => x"87e9c248",
   958 => x"48ddf2c2",
   959 => x"c27e50c0",
   960 => x"49bfccf2",
   961 => x"bffce9c2",
   962 => x"04aa714a",
   963 => x"cf87f4fb",
   964 => x"f8ffffff",
   965 => x"f0f6c24c",
   966 => x"c8c005bf",
   967 => x"c8f2c287",
   968 => x"fac102bf",
   969 => x"f8e9c287",
   970 => x"f5e649bf",
   971 => x"fce9c287",
   972 => x"48a6c458",
   973 => x"bff8e9c2",
   974 => x"c8f2c278",
   975 => x"dbc002bf",
   976 => x"4966c487",
   977 => x"a9749974",
   978 => x"87c8c002",
   979 => x"c048a6c8",
   980 => x"87e7c078",
   981 => x"c148a6c8",
   982 => x"87dfc078",
   983 => x"cf4966c4",
   984 => x"a999f8ff",
   985 => x"87c8c002",
   986 => x"c048a6cc",
   987 => x"87c5c078",
   988 => x"c148a6cc",
   989 => x"48a6c878",
   990 => x"c87866cc",
   991 => x"dec00566",
   992 => x"4966c487",
   993 => x"f2c289c2",
   994 => x"c291bfc0",
   995 => x"48bfdcf6",
   996 => x"e9c28071",
   997 => x"e9c258f8",
   998 => x"78c048fc",
   999 => x"c087d4f9",
  1000 => x"ffffcf48",
  1001 => x"f04cf8ff",
  1002 => x"264d268e",
  1003 => x"264b264c",
  1004 => x"0000004f",
  1005 => x"00000000",
  1006 => x"ffffffff",
  1007 => x"00000fc4",
  1008 => x"00000fd0",
  1009 => x"33544146",
  1010 => x"20202032",
  1011 => x"00000000",
  1012 => x"31544146",
  1013 => x"20202036",
  1014 => x"d4ff1e00",
  1015 => x"78ffc348",
  1016 => x"4f264868",
  1017 => x"48d4ff1e",
  1018 => x"ff78ffc3",
  1019 => x"e1c048d0",
  1020 => x"48d4ff78",
  1021 => x"4f2678d4",
  1022 => x"48d0ff1e",
  1023 => x"2678e0c0",
  1024 => x"d4ff1e4f",
  1025 => x"99497087",
  1026 => x"c087c602",
  1027 => x"f105a9fb",
  1028 => x"26487187",
  1029 => x"5b5e0e4f",
  1030 => x"4b710e5c",
  1031 => x"f8fe4cc0",
  1032 => x"99497087",
  1033 => x"87f9c002",
  1034 => x"02a9ecc0",
  1035 => x"c087f2c0",
  1036 => x"c002a9fb",
  1037 => x"66cc87eb",
  1038 => x"c703acb7",
  1039 => x"0266d087",
  1040 => x"537187c2",
  1041 => x"c2029971",
  1042 => x"fe84c187",
  1043 => x"497087cb",
  1044 => x"87cd0299",
  1045 => x"02a9ecc0",
  1046 => x"fbc087c7",
  1047 => x"d5ff05a9",
  1048 => x"0266d087",
  1049 => x"97c087c3",
  1050 => x"a9ecc07b",
  1051 => x"7487c405",
  1052 => x"7487c54a",
  1053 => x"8a0ac04a",
  1054 => x"4c264872",
  1055 => x"4f264b26",
  1056 => x"87d5fd1e",
  1057 => x"c04a4970",
  1058 => x"c904aaf0",
  1059 => x"aaf9c087",
  1060 => x"c087c301",
  1061 => x"c1c18af0",
  1062 => x"87c904aa",
  1063 => x"01aadac1",
  1064 => x"f7c087c3",
  1065 => x"2648728a",
  1066 => x"5b5e0e4f",
  1067 => x"f80e5d5c",
  1068 => x"c04c7186",
  1069 => x"87ecfc7e",
  1070 => x"c5c14bc0",
  1071 => x"49bf97c8",
  1072 => x"cf04a9c0",
  1073 => x"87f9fc87",
  1074 => x"c5c183c1",
  1075 => x"49bf97c8",
  1076 => x"87f106ab",
  1077 => x"97c8c5c1",
  1078 => x"87cf02bf",
  1079 => x"7087fafb",
  1080 => x"c6029949",
  1081 => x"a9ecc087",
  1082 => x"c087f105",
  1083 => x"87e9fb4b",
  1084 => x"e4fb4d70",
  1085 => x"58a6c887",
  1086 => x"7087defb",
  1087 => x"c883c14a",
  1088 => x"699749a4",
  1089 => x"da05ad49",
  1090 => x"49a4c987",
  1091 => x"c4496997",
  1092 => x"ce05a966",
  1093 => x"49a4ca87",
  1094 => x"aa496997",
  1095 => x"c187c405",
  1096 => x"c087d07e",
  1097 => x"c602adec",
  1098 => x"adfbc087",
  1099 => x"c087c405",
  1100 => x"6e7ec14b",
  1101 => x"87f5fe02",
  1102 => x"7387fdfa",
  1103 => x"268ef848",
  1104 => x"264c264d",
  1105 => x"004f264b",
  1106 => x"1e731e00",
  1107 => x"c84bd4ff",
  1108 => x"d0ff4a66",
  1109 => x"78c5c848",
  1110 => x"c148d4ff",
  1111 => x"7b1178d4",
  1112 => x"f9058ac1",
  1113 => x"48d0ff87",
  1114 => x"4b2678c4",
  1115 => x"5e0e4f26",
  1116 => x"0e5d5c5b",
  1117 => x"7e7186f8",
  1118 => x"f7c21e6e",
  1119 => x"dfff49c0",
  1120 => x"86c487d7",
  1121 => x"c4029870",
  1122 => x"f4c187e4",
  1123 => x"6e4cbfd0",
  1124 => x"87d5fc49",
  1125 => x"7058a6c8",
  1126 => x"87c50598",
  1127 => x"c148a6c4",
  1128 => x"48d0ff78",
  1129 => x"d4ff78c5",
  1130 => x"78d5c148",
  1131 => x"c14966c4",
  1132 => x"c131c689",
  1133 => x"bf97c8f4",
  1134 => x"b071484a",
  1135 => x"7808d4ff",
  1136 => x"c448d0ff",
  1137 => x"fcf6c278",
  1138 => x"d049bf97",
  1139 => x"87dd0299",
  1140 => x"d4ff78c5",
  1141 => x"78d6c148",
  1142 => x"d4ff4ac0",
  1143 => x"78ffc348",
  1144 => x"e0c082c1",
  1145 => x"87f204aa",
  1146 => x"c448d0ff",
  1147 => x"48d4ff78",
  1148 => x"ff78ffc3",
  1149 => x"78c548d0",
  1150 => x"c148d4ff",
  1151 => x"78c178d3",
  1152 => x"c448d0ff",
  1153 => x"acb7c078",
  1154 => x"87cbc206",
  1155 => x"bfc8f7c2",
  1156 => x"7e748c4b",
  1157 => x"c1029b73",
  1158 => x"c0c887dd",
  1159 => x"b7c08b4d",
  1160 => x"87c603ab",
  1161 => x"4da3c0c8",
  1162 => x"f6c24bc0",
  1163 => x"49bf97fc",
  1164 => x"cf0299d0",
  1165 => x"c21ec087",
  1166 => x"e249c0f7",
  1167 => x"86c487d9",
  1168 => x"87d84c70",
  1169 => x"1ec0eac2",
  1170 => x"49c0f7c2",
  1171 => x"7087c8e2",
  1172 => x"c21e754c",
  1173 => x"fb49c0ea",
  1174 => x"86c887ef",
  1175 => x"c5059c74",
  1176 => x"c148c087",
  1177 => x"1ec187ca",
  1178 => x"49c0f7c2",
  1179 => x"c487cde0",
  1180 => x"059b7386",
  1181 => x"6e87e3fe",
  1182 => x"acb7c04c",
  1183 => x"c287d106",
  1184 => x"c048c0f7",
  1185 => x"c080d078",
  1186 => x"c280f478",
  1187 => x"78bfccf7",
  1188 => x"01acb7c0",
  1189 => x"ff87f5fd",
  1190 => x"78c548d0",
  1191 => x"c148d4ff",
  1192 => x"78c078d3",
  1193 => x"c448d0ff",
  1194 => x"c048c178",
  1195 => x"48c087c2",
  1196 => x"4d268ef8",
  1197 => x"4b264c26",
  1198 => x"5e0e4f26",
  1199 => x"0e5d5c5b",
  1200 => x"4d7186fc",
  1201 => x"ad4c4bc0",
  1202 => x"87e8c004",
  1203 => x"1ee9c2c1",
  1204 => x"c4029c74",
  1205 => x"c24ac087",
  1206 => x"724ac187",
  1207 => x"87ddeb49",
  1208 => x"7e7086c4",
  1209 => x"056e83c1",
  1210 => x"4b7587c2",
  1211 => x"ab7584c1",
  1212 => x"87d8ff06",
  1213 => x"8efc486e",
  1214 => x"4c264d26",
  1215 => x"4f264b26",
  1216 => x"5c5b5e0e",
  1217 => x"cc4b710e",
  1218 => x"87d80266",
  1219 => x"8cf0c04c",
  1220 => x"7487d802",
  1221 => x"028ac14a",
  1222 => x"028a87d1",
  1223 => x"028a87cd",
  1224 => x"87d987c9",
  1225 => x"c5f94973",
  1226 => x"7487d287",
  1227 => x"c149c01e",
  1228 => x"7487fdd9",
  1229 => x"c149731e",
  1230 => x"c887f5d9",
  1231 => x"264c2686",
  1232 => x"0e4f264b",
  1233 => x"5d5c5b5e",
  1234 => x"7186fc0e",
  1235 => x"91de494c",
  1236 => x"4de0f8c2",
  1237 => x"6d978571",
  1238 => x"87dcc102",
  1239 => x"bfd0f8c2",
  1240 => x"71817449",
  1241 => x"7087d3fd",
  1242 => x"0298487e",
  1243 => x"c287f2c0",
  1244 => x"704bd4f8",
  1245 => x"fe49cb4a",
  1246 => x"7487e9f6",
  1247 => x"c193cc4b",
  1248 => x"c483d4f4",
  1249 => x"c4cfc183",
  1250 => x"c149747b",
  1251 => x"7587e9c4",
  1252 => x"ccf4c17b",
  1253 => x"1e49bf97",
  1254 => x"49d4f8c2",
  1255 => x"c487e1fd",
  1256 => x"c1497486",
  1257 => x"c087d1c4",
  1258 => x"ecc5c149",
  1259 => x"f8f6c287",
  1260 => x"4950c048",
  1261 => x"87cbe2c0",
  1262 => x"4d268efc",
  1263 => x"4b264c26",
  1264 => x"00004f26",
  1265 => x"64616f4c",
  1266 => x"2e676e69",
  1267 => x"1e002e2e",
  1268 => x"4b711e73",
  1269 => x"d0f8c249",
  1270 => x"fb7181bf",
  1271 => x"4a7087dc",
  1272 => x"87c4029a",
  1273 => x"87dbe649",
  1274 => x"48d0f8c2",
  1275 => x"497378c0",
  1276 => x"2687fac1",
  1277 => x"1e4f264b",
  1278 => x"4b711e73",
  1279 => x"024aa3c4",
  1280 => x"c187d0c1",
  1281 => x"87dc028a",
  1282 => x"f2c0028a",
  1283 => x"c1058a87",
  1284 => x"f8c287d3",
  1285 => x"c102bfd0",
  1286 => x"c14887cb",
  1287 => x"d4f8c288",
  1288 => x"87c1c158",
  1289 => x"bfd0f8c2",
  1290 => x"c289c649",
  1291 => x"c059d4f8",
  1292 => x"c003a9b7",
  1293 => x"f8c287ef",
  1294 => x"78c048d0",
  1295 => x"c287e6c0",
  1296 => x"02bfccf8",
  1297 => x"f8c287df",
  1298 => x"c148bfd0",
  1299 => x"d4f8c280",
  1300 => x"c287d258",
  1301 => x"02bfccf8",
  1302 => x"f8c287cb",
  1303 => x"c648bfd0",
  1304 => x"d4f8c280",
  1305 => x"c4497358",
  1306 => x"264b2687",
  1307 => x"5b5e0e4f",
  1308 => x"f00e5d5c",
  1309 => x"59a6d086",
  1310 => x"4dc0eac2",
  1311 => x"f8c24cc0",
  1312 => x"78c148cc",
  1313 => x"c048a6c8",
  1314 => x"c27e7578",
  1315 => x"48bfd0f8",
  1316 => x"c106a8c0",
  1317 => x"a6c887c0",
  1318 => x"c27e755c",
  1319 => x"9848c0ea",
  1320 => x"87f2c002",
  1321 => x"c14d66c4",
  1322 => x"cc1ee9c2",
  1323 => x"87c40266",
  1324 => x"87c24cc0",
  1325 => x"49744cc1",
  1326 => x"c487c2e4",
  1327 => x"c17e7086",
  1328 => x"4866c885",
  1329 => x"a6cc80c1",
  1330 => x"d0f8c258",
  1331 => x"c503adbf",
  1332 => x"ff056e87",
  1333 => x"4d6e87d1",
  1334 => x"9d754cc0",
  1335 => x"87dcc302",
  1336 => x"1ee9c2c1",
  1337 => x"c70266cc",
  1338 => x"48a6c887",
  1339 => x"87c578c0",
  1340 => x"c148a6c8",
  1341 => x"4966c878",
  1342 => x"c487c2e3",
  1343 => x"487e7086",
  1344 => x"e4c20298",
  1345 => x"81cb4987",
  1346 => x"d0496997",
  1347 => x"d4c10299",
  1348 => x"cc497487",
  1349 => x"d4f4c191",
  1350 => x"cfcfc181",
  1351 => x"c381c879",
  1352 => x"497451ff",
  1353 => x"f8c291de",
  1354 => x"85714de0",
  1355 => x"7d97c1c2",
  1356 => x"c049a5c1",
  1357 => x"f2c251e0",
  1358 => x"02bf97d0",
  1359 => x"84c187d2",
  1360 => x"c24ba5c2",
  1361 => x"db4ad0f2",
  1362 => x"d7effe49",
  1363 => x"87d9c187",
  1364 => x"c049a5cd",
  1365 => x"c284c151",
  1366 => x"4a6e4ba5",
  1367 => x"effe49cb",
  1368 => x"c4c187c2",
  1369 => x"cc497487",
  1370 => x"d4f4c191",
  1371 => x"c3cdc181",
  1372 => x"d0f2c279",
  1373 => x"d802bf97",
  1374 => x"de497487",
  1375 => x"c284c191",
  1376 => x"714be0f8",
  1377 => x"d0f2c283",
  1378 => x"fe49dd4a",
  1379 => x"d887d5ee",
  1380 => x"de4b7487",
  1381 => x"e0f8c293",
  1382 => x"49a3cb83",
  1383 => x"84c151c0",
  1384 => x"cb4a6e73",
  1385 => x"fbedfe49",
  1386 => x"4866c887",
  1387 => x"a6cc80c1",
  1388 => x"03acc758",
  1389 => x"6e87c5c0",
  1390 => x"87e4fc05",
  1391 => x"c003acc7",
  1392 => x"f8c287e4",
  1393 => x"78c048cc",
  1394 => x"91cc4974",
  1395 => x"81d4f4c1",
  1396 => x"79c3cdc1",
  1397 => x"91de4974",
  1398 => x"81e0f8c2",
  1399 => x"84c151c0",
  1400 => x"ff04acc7",
  1401 => x"f5c187dc",
  1402 => x"50c048f0",
  1403 => x"d9c180f7",
  1404 => x"d8c140dd",
  1405 => x"80c878d0",
  1406 => x"78f7cfc1",
  1407 => x"c04966cc",
  1408 => x"f087f5fa",
  1409 => x"264d268e",
  1410 => x"264b264c",
  1411 => x"0000004f",
  1412 => x"61422080",
  1413 => x"1e006b63",
  1414 => x"4b711e73",
  1415 => x"c191cc49",
  1416 => x"c881d4f4",
  1417 => x"f4c14aa1",
  1418 => x"501248c8",
  1419 => x"c14aa1c9",
  1420 => x"1248c8c5",
  1421 => x"c181ca50",
  1422 => x"1148ccf4",
  1423 => x"ccf4c150",
  1424 => x"1e49bf97",
  1425 => x"f7f249c0",
  1426 => x"f8497387",
  1427 => x"8efc87df",
  1428 => x"4f264b26",
  1429 => x"c049c01e",
  1430 => x"2687fefa",
  1431 => x"4a711e4f",
  1432 => x"c191cc49",
  1433 => x"c881d4f4",
  1434 => x"f8f6c281",
  1435 => x"c0501148",
  1436 => x"fe49a2f0",
  1437 => x"c087d5e8",
  1438 => x"87c7d749",
  1439 => x"ff1e4f26",
  1440 => x"ffc34ad4",
  1441 => x"48d0ff7a",
  1442 => x"de78e1c0",
  1443 => x"487a717a",
  1444 => x"7028b7c8",
  1445 => x"d048717a",
  1446 => x"7a7028b7",
  1447 => x"b7d84871",
  1448 => x"ff7a7028",
  1449 => x"e0c048d0",
  1450 => x"0e4f2678",
  1451 => x"5d5c5b5e",
  1452 => x"7186f40e",
  1453 => x"91cc494d",
  1454 => x"81d4f4c1",
  1455 => x"ca4aa1c8",
  1456 => x"a6c47ea1",
  1457 => x"f4f6c248",
  1458 => x"976e78bf",
  1459 => x"66c44bbf",
  1460 => x"122c734c",
  1461 => x"58a6cc48",
  1462 => x"84c19c70",
  1463 => x"699781c9",
  1464 => x"04acb749",
  1465 => x"4cc087c2",
  1466 => x"4abf976e",
  1467 => x"724966c8",
  1468 => x"c4b9ff31",
  1469 => x"48749966",
  1470 => x"4a703072",
  1471 => x"f8f6c2b1",
  1472 => x"f9fd7159",
  1473 => x"c21ec787",
  1474 => x"1ebfc8f8",
  1475 => x"1ed4f4c1",
  1476 => x"97f8f6c2",
  1477 => x"f4c149bf",
  1478 => x"c0497587",
  1479 => x"e887d9f6",
  1480 => x"264d268e",
  1481 => x"264b264c",
  1482 => x"1e731e4f",
  1483 => x"fd494b71",
  1484 => x"497387f9",
  1485 => x"2687f4fd",
  1486 => x"1e4f264b",
  1487 => x"4b711e73",
  1488 => x"024aa3c2",
  1489 => x"8ac187d6",
  1490 => x"87e2c005",
  1491 => x"bfc8f8c2",
  1492 => x"4887db02",
  1493 => x"f8c288c1",
  1494 => x"87d258cc",
  1495 => x"bfccf8c2",
  1496 => x"c287cb02",
  1497 => x"48bfc8f8",
  1498 => x"f8c280c1",
  1499 => x"1ec758cc",
  1500 => x"bfc8f8c2",
  1501 => x"d4f4c11e",
  1502 => x"f8f6c21e",
  1503 => x"cc49bf97",
  1504 => x"c0497387",
  1505 => x"f487f1f4",
  1506 => x"264b268e",
  1507 => x"5b5e0e4f",
  1508 => x"ff0e5d5c",
  1509 => x"e4c086cc",
  1510 => x"a6cc59a6",
  1511 => x"c478c048",
  1512 => x"c478c080",
  1513 => x"66c8c180",
  1514 => x"c180c478",
  1515 => x"c180c478",
  1516 => x"ccf8c278",
  1517 => x"e078c148",
  1518 => x"c4e187ea",
  1519 => x"87d9e087",
  1520 => x"fbc04c70",
  1521 => x"f3c102ac",
  1522 => x"66e0c087",
  1523 => x"87e8c105",
  1524 => x"4a66c4c1",
  1525 => x"7e6a82c4",
  1526 => x"48e4f0c1",
  1527 => x"4120496e",
  1528 => x"51104120",
  1529 => x"4866c4c1",
  1530 => x"78d7d8c1",
  1531 => x"81c7496a",
  1532 => x"c4c15174",
  1533 => x"81c84966",
  1534 => x"a6d851c1",
  1535 => x"c178c248",
  1536 => x"c94966c4",
  1537 => x"c151c081",
  1538 => x"ca4966c4",
  1539 => x"c151c081",
  1540 => x"6a1ed81e",
  1541 => x"ff81c849",
  1542 => x"c887fadf",
  1543 => x"66c8c186",
  1544 => x"01a8c048",
  1545 => x"a6d087c7",
  1546 => x"cf78c148",
  1547 => x"66c8c187",
  1548 => x"d888c148",
  1549 => x"87c458a6",
  1550 => x"87c5dfff",
  1551 => x"cd029c74",
  1552 => x"66d087da",
  1553 => x"66ccc148",
  1554 => x"cfcd03a8",
  1555 => x"48a6c887",
  1556 => x"ff7e78c0",
  1557 => x"7087c2de",
  1558 => x"acd0c14c",
  1559 => x"87e7c205",
  1560 => x"6e48a6c4",
  1561 => x"87d8e078",
  1562 => x"cc487e70",
  1563 => x"c506a866",
  1564 => x"48a6cc87",
  1565 => x"ddff786e",
  1566 => x"4c7087df",
  1567 => x"05acecc0",
  1568 => x"d087eec1",
  1569 => x"91cc4966",
  1570 => x"8166c4c1",
  1571 => x"6a4aa1c4",
  1572 => x"4aa1c84d",
  1573 => x"d9c1526e",
  1574 => x"dcff79dd",
  1575 => x"4c7087fb",
  1576 => x"87d9029c",
  1577 => x"02acfbc0",
  1578 => x"557487d3",
  1579 => x"87e9dcff",
  1580 => x"029c4c70",
  1581 => x"fbc087c7",
  1582 => x"edff05ac",
  1583 => x"55e0c087",
  1584 => x"c055c1c2",
  1585 => x"e0c07d97",
  1586 => x"66c44866",
  1587 => x"87db05a8",
  1588 => x"d44866d0",
  1589 => x"ca04a866",
  1590 => x"4866d087",
  1591 => x"a6d480c1",
  1592 => x"d487c858",
  1593 => x"88c14866",
  1594 => x"ff58a6d8",
  1595 => x"7087eadb",
  1596 => x"acd0c14c",
  1597 => x"dc87c905",
  1598 => x"80c14866",
  1599 => x"58a6e0c0",
  1600 => x"02acd0c1",
  1601 => x"6e87d9fd",
  1602 => x"66e0c048",
  1603 => x"ebc905a8",
  1604 => x"a6e4c087",
  1605 => x"7478c048",
  1606 => x"88fbc048",
  1607 => x"7058a6c8",
  1608 => x"ddc90298",
  1609 => x"88cb4887",
  1610 => x"7058a6c8",
  1611 => x"cfc10298",
  1612 => x"88c94887",
  1613 => x"7058a6c8",
  1614 => x"ffc30298",
  1615 => x"88c44887",
  1616 => x"7058a6c8",
  1617 => x"87cf0298",
  1618 => x"c888c148",
  1619 => x"987058a6",
  1620 => x"87e8c302",
  1621 => x"c887dcc8",
  1622 => x"f0c048a6",
  1623 => x"f8d9ff78",
  1624 => x"c04c7087",
  1625 => x"c002acec",
  1626 => x"a6cc87c3",
  1627 => x"acecc05c",
  1628 => x"ff87cd02",
  1629 => x"7087e2d9",
  1630 => x"acecc04c",
  1631 => x"87f3ff05",
  1632 => x"02acecc0",
  1633 => x"ff87c4c0",
  1634 => x"c087ced9",
  1635 => x"d81eca1e",
  1636 => x"91cc4966",
  1637 => x"4866ccc1",
  1638 => x"a6cc8071",
  1639 => x"4866c858",
  1640 => x"a6d080c4",
  1641 => x"bf66cc58",
  1642 => x"e8d9ff49",
  1643 => x"de1ec187",
  1644 => x"bf66d41e",
  1645 => x"dcd9ff49",
  1646 => x"7086d087",
  1647 => x"08c04849",
  1648 => x"a6ecc088",
  1649 => x"06a8c058",
  1650 => x"c087eec0",
  1651 => x"dd4866e8",
  1652 => x"e4c003a8",
  1653 => x"bf66c487",
  1654 => x"66e8c049",
  1655 => x"51e0c081",
  1656 => x"4966e8c0",
  1657 => x"66c481c1",
  1658 => x"c1c281bf",
  1659 => x"66e8c051",
  1660 => x"c481c249",
  1661 => x"c081bf66",
  1662 => x"c1486e51",
  1663 => x"6e78d7d8",
  1664 => x"d881c849",
  1665 => x"496e5166",
  1666 => x"66dc81c9",
  1667 => x"ca496e51",
  1668 => x"5166c881",
  1669 => x"c14866d8",
  1670 => x"58a6dc80",
  1671 => x"d44866d0",
  1672 => x"c004a866",
  1673 => x"66d087cb",
  1674 => x"d480c148",
  1675 => x"d1c558a6",
  1676 => x"4866d487",
  1677 => x"a6d888c1",
  1678 => x"87c6c558",
  1679 => x"87c0d9ff",
  1680 => x"58a6ecc0",
  1681 => x"87f8d8ff",
  1682 => x"58a6f0c0",
  1683 => x"05a8ecc0",
  1684 => x"a687c9c0",
  1685 => x"66e8c048",
  1686 => x"87c4c078",
  1687 => x"87f9d5ff",
  1688 => x"cc4966d0",
  1689 => x"66c4c191",
  1690 => x"c8807148",
  1691 => x"66c458a6",
  1692 => x"c482c84a",
  1693 => x"81ca4966",
  1694 => x"5166e8c0",
  1695 => x"4966ecc0",
  1696 => x"e8c081c1",
  1697 => x"48c18966",
  1698 => x"49703071",
  1699 => x"977189c1",
  1700 => x"f4f6c27a",
  1701 => x"e8c049bf",
  1702 => x"6a972966",
  1703 => x"9871484a",
  1704 => x"58a6f4c0",
  1705 => x"c44866c4",
  1706 => x"58a6cc80",
  1707 => x"4dbf66c8",
  1708 => x"4866e0c0",
  1709 => x"c002a86e",
  1710 => x"7ec087c5",
  1711 => x"c187c2c0",
  1712 => x"c01e6e7e",
  1713 => x"49751ee0",
  1714 => x"87c9d5ff",
  1715 => x"4c7086c8",
  1716 => x"06acb7c0",
  1717 => x"7487d4c1",
  1718 => x"bf66c885",
  1719 => x"81e0c049",
  1720 => x"c14b8975",
  1721 => x"714af0f0",
  1722 => x"87f8d8fe",
  1723 => x"7e7585c2",
  1724 => x"4866e4c0",
  1725 => x"e8c080c1",
  1726 => x"f0c058a6",
  1727 => x"81c14966",
  1728 => x"c002a970",
  1729 => x"4dc087c5",
  1730 => x"c187c2c0",
  1731 => x"cc1e754d",
  1732 => x"c049bf66",
  1733 => x"66c481e0",
  1734 => x"c81e7189",
  1735 => x"d3ff4966",
  1736 => x"86c887f3",
  1737 => x"01a8b7c0",
  1738 => x"c087c5ff",
  1739 => x"c00266e4",
  1740 => x"66c487d3",
  1741 => x"c081c949",
  1742 => x"c45166e4",
  1743 => x"dac14866",
  1744 => x"cec078eb",
  1745 => x"4966c487",
  1746 => x"51c281c9",
  1747 => x"c14866c4",
  1748 => x"d078e9dc",
  1749 => x"66d44866",
  1750 => x"cbc004a8",
  1751 => x"4866d087",
  1752 => x"a6d480c1",
  1753 => x"87dac058",
  1754 => x"c14866d4",
  1755 => x"58a6d888",
  1756 => x"ff87cfc0",
  1757 => x"7087cad2",
  1758 => x"87c6c04c",
  1759 => x"87c1d2ff",
  1760 => x"66dc4c70",
  1761 => x"c080c148",
  1762 => x"7458a6e0",
  1763 => x"cbc0029c",
  1764 => x"4866d087",
  1765 => x"a866ccc1",
  1766 => x"87f1f204",
  1767 => x"c74866d0",
  1768 => x"e1c003a8",
  1769 => x"4c66d087",
  1770 => x"48ccf8c2",
  1771 => x"497478c0",
  1772 => x"c4c191cc",
  1773 => x"a1c48166",
  1774 => x"c04a6a4a",
  1775 => x"84c17952",
  1776 => x"ff04acc7",
  1777 => x"e0c087e2",
  1778 => x"e2c00266",
  1779 => x"66c4c187",
  1780 => x"81d4c149",
  1781 => x"4a66c4c1",
  1782 => x"c082dcc1",
  1783 => x"ddd9c152",
  1784 => x"66c4c179",
  1785 => x"81d8c149",
  1786 => x"79f4f0c1",
  1787 => x"c187d6c0",
  1788 => x"c14966c4",
  1789 => x"c4c181d4",
  1790 => x"d8c14a66",
  1791 => x"fcf0c182",
  1792 => x"d4d9c17a",
  1793 => x"66c4c179",
  1794 => x"81e0c149",
  1795 => x"79fbdcc1",
  1796 => x"87e4cfff",
  1797 => x"ff4866cc",
  1798 => x"4d268ecc",
  1799 => x"4b264c26",
  1800 => x"00004f26",
  1801 => x"64616f4c",
  1802 => x"202e2a20",
  1803 => x"00000000",
  1804 => x"0000203a",
  1805 => x"61422080",
  1806 => x"00006b63",
  1807 => x"78452080",
  1808 => x"1e007469",
  1809 => x"f8c21ec7",
  1810 => x"c11ebfc8",
  1811 => x"c21ed4f4",
  1812 => x"bf97f8f6",
  1813 => x"87f5ec49",
  1814 => x"49d4f4c1",
  1815 => x"87e6e2c0",
  1816 => x"4f268ef4",
  1817 => x"c81e731e",
  1818 => x"f8c287c3",
  1819 => x"50c048d4",
  1820 => x"48ecf5c1",
  1821 => x"78f4f3c1",
  1822 => x"49a0e8fe",
  1823 => x"87c6e2c0",
  1824 => x"e0c049c7",
  1825 => x"49c187f2",
  1826 => x"87cde2c0",
  1827 => x"c348d4ff",
  1828 => x"ddfe78ff",
  1829 => x"987087da",
  1830 => x"fe87cd02",
  1831 => x"7087d6e7",
  1832 => x"87c40298",
  1833 => x"87c24ac1",
  1834 => x"9a724ac0",
  1835 => x"c187c802",
  1836 => x"fe49c0f4",
  1837 => x"c287f0cf",
  1838 => x"c048c8f8",
  1839 => x"f8f6c278",
  1840 => x"4950c048",
  1841 => x"c087fcfd",
  1842 => x"7087eaf5",
  1843 => x"cb029b4b",
  1844 => x"f0f5c187",
  1845 => x"df49c75b",
  1846 => x"87c687de",
  1847 => x"e0c049c0",
  1848 => x"c2c387f7",
  1849 => x"d8e2c087",
  1850 => x"ecefc087",
  1851 => x"87f5ff87",
  1852 => x"4f264b26",
  1853 => x"746f6f42",
  1854 => x"2e676e69",
  1855 => x"00002e2e",
  1856 => x"4f204453",
  1857 => x"0000004b",
  1858 => x"00000000",
  1859 => x"00000000",
  1860 => x"00000001",
  1861 => x"00001343",
  1862 => x"00002e20",
  1863 => x"00000000",
  1864 => x"00001343",
  1865 => x"00002e3e",
  1866 => x"00000000",
  1867 => x"00001343",
  1868 => x"00002e5c",
  1869 => x"00000000",
  1870 => x"00001343",
  1871 => x"00002e7a",
  1872 => x"00000000",
  1873 => x"00001343",
  1874 => x"00002e98",
  1875 => x"00000000",
  1876 => x"00001343",
  1877 => x"00002eb6",
  1878 => x"00000000",
  1879 => x"00001343",
  1880 => x"00002ed4",
  1881 => x"00000000",
  1882 => x"0000165d",
  1883 => x"00000000",
  1884 => x"00000000",
  1885 => x"000013f7",
  1886 => x"00000000",
  1887 => x"00000000",
  1888 => x"db86fc1e",
  1889 => x"fc7e7087",
  1890 => x"1e4f268e",
  1891 => x"c048f0fe",
  1892 => x"7909cd78",
  1893 => x"1e4f2609",
  1894 => x"49c0f6c1",
  1895 => x"4f2687ed",
  1896 => x"bff0fe1e",
  1897 => x"1e4f2648",
  1898 => x"c148f0fe",
  1899 => x"1e4f2678",
  1900 => x"c048f0fe",
  1901 => x"1e4f2678",
  1902 => x"52c04a71",
  1903 => x"0e4f2651",
  1904 => x"5d5c5b5e",
  1905 => x"7186f40e",
  1906 => x"7e6d974d",
  1907 => x"974ca5c1",
  1908 => x"a6c8486c",
  1909 => x"c4486e58",
  1910 => x"c505a866",
  1911 => x"c048ff87",
  1912 => x"caff87e6",
  1913 => x"49a5c287",
  1914 => x"714b6c97",
  1915 => x"6b974ba3",
  1916 => x"7e6c974b",
  1917 => x"80c1486e",
  1918 => x"c758a6c8",
  1919 => x"58a6cc98",
  1920 => x"fe7c9770",
  1921 => x"487387e1",
  1922 => x"4d268ef4",
  1923 => x"4b264c26",
  1924 => x"5e0e4f26",
  1925 => x"f40e5c5b",
  1926 => x"d84c7186",
  1927 => x"ffc34a66",
  1928 => x"4ba4c29a",
  1929 => x"73496c97",
  1930 => x"517249a1",
  1931 => x"6e7e6c97",
  1932 => x"c880c148",
  1933 => x"98c758a6",
  1934 => x"7058a6cc",
  1935 => x"268ef454",
  1936 => x"264b264c",
  1937 => x"86fc1e4f",
  1938 => x"e087e4fd",
  1939 => x"c0494abf",
  1940 => x"0299c0e0",
  1941 => x"1e7287cb",
  1942 => x"49f4fbc2",
  1943 => x"c487f3fe",
  1944 => x"87fcfc86",
  1945 => x"fefc7e70",
  1946 => x"268efc87",
  1947 => x"fbc21e4f",
  1948 => x"c2fd49f4",
  1949 => x"c5f9c187",
  1950 => x"87cffc49",
  1951 => x"2687edc3",
  1952 => x"5b5e0e4f",
  1953 => x"fc0e5d5c",
  1954 => x"ff7e7186",
  1955 => x"fbc24dd4",
  1956 => x"eafc49f4",
  1957 => x"c04b7087",
  1958 => x"c204abb7",
  1959 => x"f0c387f8",
  1960 => x"87c905ab",
  1961 => x"48e4fdc1",
  1962 => x"d9c278c1",
  1963 => x"abe0c387",
  1964 => x"c187c905",
  1965 => x"c148e8fd",
  1966 => x"87cac278",
  1967 => x"bfe8fdc1",
  1968 => x"c287c602",
  1969 => x"c24ca3c0",
  1970 => x"c14c7387",
  1971 => x"02bfe4fd",
  1972 => x"7487e0c0",
  1973 => x"29b7c449",
  1974 => x"c0ffc191",
  1975 => x"cf4a7481",
  1976 => x"c192c29a",
  1977 => x"70307248",
  1978 => x"72baff4a",
  1979 => x"70986948",
  1980 => x"7487db79",
  1981 => x"29b7c449",
  1982 => x"c0ffc191",
  1983 => x"cf4a7481",
  1984 => x"c392c29a",
  1985 => x"70307248",
  1986 => x"b069484a",
  1987 => x"056e7970",
  1988 => x"ff87e7c0",
  1989 => x"e1c848d0",
  1990 => x"c17dc578",
  1991 => x"02bfe8fd",
  1992 => x"e0c387c3",
  1993 => x"e4fdc17d",
  1994 => x"87c302bf",
  1995 => x"737df0c3",
  1996 => x"48d0ff7d",
  1997 => x"c078e1c8",
  1998 => x"fdc178e0",
  1999 => x"78c048e8",
  2000 => x"48e4fdc1",
  2001 => x"fbc278c0",
  2002 => x"f2f949f4",
  2003 => x"c04b7087",
  2004 => x"fd03abb7",
  2005 => x"48c087c8",
  2006 => x"4d268efc",
  2007 => x"4b264c26",
  2008 => x"00004f26",
  2009 => x"00000000",
  2010 => x"00000000",
  2011 => x"724ac01e",
  2012 => x"c191c449",
  2013 => x"c081c0ff",
  2014 => x"d082c179",
  2015 => x"ee04aab7",
  2016 => x"0e4f2687",
  2017 => x"5d5c5b5e",
  2018 => x"f84d710e",
  2019 => x"4a7587e1",
  2020 => x"922ab7c4",
  2021 => x"82c0ffc1",
  2022 => x"9ccf4c75",
  2023 => x"496a94c2",
  2024 => x"c32b744b",
  2025 => x"7448c29b",
  2026 => x"ff4c7030",
  2027 => x"714874bc",
  2028 => x"f77a7098",
  2029 => x"487387f1",
  2030 => x"4c264d26",
  2031 => x"4f264b26",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"00000000",
  2035 => x"00000000",
  2036 => x"00000000",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00000000",
  2040 => x"00000000",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00000000",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"00000000",
  2048 => x"48d0ff1e",
  2049 => x"7178e1c8",
  2050 => x"08d4ff48",
  2051 => x"1e4f2678",
  2052 => x"c848d0ff",
  2053 => x"487178e1",
  2054 => x"7808d4ff",
  2055 => x"ff4866c4",
  2056 => x"267808d4",
  2057 => x"4a711e4f",
  2058 => x"1e4966c4",
  2059 => x"deff4972",
  2060 => x"48d0ff87",
  2061 => x"fc78e0c0",
  2062 => x"1e4f268e",
  2063 => x"4a711e73",
  2064 => x"abb7c24b",
  2065 => x"a387c803",
  2066 => x"ffc34a49",
  2067 => x"ce87c79a",
  2068 => x"c34a49a3",
  2069 => x"66c89aff",
  2070 => x"49721e49",
  2071 => x"fc87c6ff",
  2072 => x"264b268e",
  2073 => x"d0ff1e4f",
  2074 => x"78c9c848",
  2075 => x"d4ff4871",
  2076 => x"4f267808",
  2077 => x"494a711e",
  2078 => x"d0ff87eb",
  2079 => x"2678c848",
  2080 => x"1e731e4f",
  2081 => x"fcc24b71",
  2082 => x"c302bfcc",
  2083 => x"87ebc287",
  2084 => x"c848d0ff",
  2085 => x"487378c9",
  2086 => x"ffb0e0c0",
  2087 => x"c27808d4",
  2088 => x"c048c0fc",
  2089 => x"0266c878",
  2090 => x"ffc387c5",
  2091 => x"c087c249",
  2092 => x"c8fcc249",
  2093 => x"0266cc59",
  2094 => x"d5c587c6",
  2095 => x"87c44ad5",
  2096 => x"4affffcf",
  2097 => x"5accfcc2",
  2098 => x"48ccfcc2",
  2099 => x"4b2678c1",
  2100 => x"5e0e4f26",
  2101 => x"0e5d5c5b",
  2102 => x"fcc24d71",
  2103 => x"754bbfc8",
  2104 => x"87cb029d",
  2105 => x"c291c849",
  2106 => x"714af8c1",
  2107 => x"c287c482",
  2108 => x"c04af8c5",
  2109 => x"7349124c",
  2110 => x"c4fcc299",
  2111 => x"b87148bf",
  2112 => x"7808d4ff",
  2113 => x"842bb7c1",
  2114 => x"04acb7c8",
  2115 => x"fcc287e7",
  2116 => x"c848bfc0",
  2117 => x"c4fcc280",
  2118 => x"264d2658",
  2119 => x"264b264c",
  2120 => x"1e731e4f",
  2121 => x"4a134b71",
  2122 => x"87cb029a",
  2123 => x"e1fe4972",
  2124 => x"9a4a1387",
  2125 => x"2687f505",
  2126 => x"1e4f264b",
  2127 => x"bfc0fcc2",
  2128 => x"c0fcc249",
  2129 => x"78a1c148",
  2130 => x"a9b7c0c4",
  2131 => x"ff87db03",
  2132 => x"fcc248d4",
  2133 => x"c278bfc4",
  2134 => x"49bfc0fc",
  2135 => x"48c0fcc2",
  2136 => x"c478a1c1",
  2137 => x"04a9b7c0",
  2138 => x"d0ff87e5",
  2139 => x"c278c848",
  2140 => x"c048ccfc",
  2141 => x"004f2678",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"5f000000",
  2145 => x"0000005f",
  2146 => x"00030300",
  2147 => x"00000303",
  2148 => x"147f7f14",
  2149 => x"00147f7f",
  2150 => x"6b2e2400",
  2151 => x"00123a6b",
  2152 => x"18366a4c",
  2153 => x"0032566c",
  2154 => x"594f7e30",
  2155 => x"40683a77",
  2156 => x"07040000",
  2157 => x"00000003",
  2158 => x"3e1c0000",
  2159 => x"00004163",
  2160 => x"63410000",
  2161 => x"00001c3e",
  2162 => x"1c3e2a08",
  2163 => x"082a3e1c",
  2164 => x"3e080800",
  2165 => x"0008083e",
  2166 => x"e0800000",
  2167 => x"00000060",
  2168 => x"08080800",
  2169 => x"00080808",
  2170 => x"60000000",
  2171 => x"00000060",
  2172 => x"18306040",
  2173 => x"0103060c",
  2174 => x"597f3e00",
  2175 => x"003e7f4d",
  2176 => x"7f060400",
  2177 => x"0000007f",
  2178 => x"71634200",
  2179 => x"00464f59",
  2180 => x"49632200",
  2181 => x"00367f49",
  2182 => x"13161c18",
  2183 => x"00107f7f",
  2184 => x"45672700",
  2185 => x"00397d45",
  2186 => x"4b7e3c00",
  2187 => x"00307949",
  2188 => x"71010100",
  2189 => x"00070f79",
  2190 => x"497f3600",
  2191 => x"00367f49",
  2192 => x"494f0600",
  2193 => x"001e3f69",
  2194 => x"66000000",
  2195 => x"00000066",
  2196 => x"e6800000",
  2197 => x"00000066",
  2198 => x"14080800",
  2199 => x"00222214",
  2200 => x"14141400",
  2201 => x"00141414",
  2202 => x"14222200",
  2203 => x"00080814",
  2204 => x"51030200",
  2205 => x"00060f59",
  2206 => x"5d417f3e",
  2207 => x"001e1f55",
  2208 => x"097f7e00",
  2209 => x"007e7f09",
  2210 => x"497f7f00",
  2211 => x"00367f49",
  2212 => x"633e1c00",
  2213 => x"00414141",
  2214 => x"417f7f00",
  2215 => x"001c3e63",
  2216 => x"497f7f00",
  2217 => x"00414149",
  2218 => x"097f7f00",
  2219 => x"00010109",
  2220 => x"417f3e00",
  2221 => x"007a7b49",
  2222 => x"087f7f00",
  2223 => x"007f7f08",
  2224 => x"7f410000",
  2225 => x"0000417f",
  2226 => x"40602000",
  2227 => x"003f7f40",
  2228 => x"1c087f7f",
  2229 => x"00416336",
  2230 => x"407f7f00",
  2231 => x"00404040",
  2232 => x"0c067f7f",
  2233 => x"007f7f06",
  2234 => x"0c067f7f",
  2235 => x"007f7f18",
  2236 => x"417f3e00",
  2237 => x"003e7f41",
  2238 => x"097f7f00",
  2239 => x"00060f09",
  2240 => x"61417f3e",
  2241 => x"00407e7f",
  2242 => x"097f7f00",
  2243 => x"00667f19",
  2244 => x"4d6f2600",
  2245 => x"00327b59",
  2246 => x"7f010100",
  2247 => x"0001017f",
  2248 => x"407f3f00",
  2249 => x"003f7f40",
  2250 => x"703f0f00",
  2251 => x"000f3f70",
  2252 => x"18307f7f",
  2253 => x"007f7f30",
  2254 => x"1c366341",
  2255 => x"4163361c",
  2256 => x"7c060301",
  2257 => x"0103067c",
  2258 => x"4d597161",
  2259 => x"00414347",
  2260 => x"7f7f0000",
  2261 => x"00004141",
  2262 => x"0c060301",
  2263 => x"40603018",
  2264 => x"41410000",
  2265 => x"00007f7f",
  2266 => x"03060c08",
  2267 => x"00080c06",
  2268 => x"80808080",
  2269 => x"00808080",
  2270 => x"03000000",
  2271 => x"00000407",
  2272 => x"54742000",
  2273 => x"00787c54",
  2274 => x"447f7f00",
  2275 => x"00387c44",
  2276 => x"447c3800",
  2277 => x"00004444",
  2278 => x"447c3800",
  2279 => x"007f7f44",
  2280 => x"547c3800",
  2281 => x"00185c54",
  2282 => x"7f7e0400",
  2283 => x"00000505",
  2284 => x"a4bc1800",
  2285 => x"007cfca4",
  2286 => x"047f7f00",
  2287 => x"00787c04",
  2288 => x"3d000000",
  2289 => x"0000407d",
  2290 => x"80808000",
  2291 => x"00007dfd",
  2292 => x"107f7f00",
  2293 => x"00446c38",
  2294 => x"3f000000",
  2295 => x"0000407f",
  2296 => x"180c7c7c",
  2297 => x"00787c0c",
  2298 => x"047c7c00",
  2299 => x"00787c04",
  2300 => x"447c3800",
  2301 => x"00387c44",
  2302 => x"24fcfc00",
  2303 => x"00183c24",
  2304 => x"243c1800",
  2305 => x"00fcfc24",
  2306 => x"047c7c00",
  2307 => x"00080c04",
  2308 => x"545c4800",
  2309 => x"00207454",
  2310 => x"7f3f0400",
  2311 => x"00004444",
  2312 => x"407c3c00",
  2313 => x"007c7c40",
  2314 => x"603c1c00",
  2315 => x"001c3c60",
  2316 => x"30607c3c",
  2317 => x"003c7c60",
  2318 => x"10386c44",
  2319 => x"00446c38",
  2320 => x"e0bc1c00",
  2321 => x"001c3c60",
  2322 => x"74644400",
  2323 => x"00444c5c",
  2324 => x"3e080800",
  2325 => x"00414177",
  2326 => x"7f000000",
  2327 => x"0000007f",
  2328 => x"77414100",
  2329 => x"0008083e",
  2330 => x"03010102",
  2331 => x"00010202",
  2332 => x"7f7f7f7f",
  2333 => x"007f7f7f",
  2334 => x"1c1c0808",
  2335 => x"7f7f3e3e",
  2336 => x"3e3e7f7f",
  2337 => x"08081c1c",
  2338 => x"7c181000",
  2339 => x"0010187c",
  2340 => x"7c301000",
  2341 => x"0010307c",
  2342 => x"60603010",
  2343 => x"00061e78",
  2344 => x"183c6642",
  2345 => x"0042663c",
  2346 => x"c26a3878",
  2347 => x"00386cc6",
  2348 => x"60000060",
  2349 => x"00600000",
  2350 => x"5c5b5e0e",
  2351 => x"86fc0e5d",
  2352 => x"fcc27e71",
  2353 => x"c04cbfd4",
  2354 => x"c41ec04b",
  2355 => x"c402ab66",
  2356 => x"c24dc087",
  2357 => x"754dc187",
  2358 => x"ee49731e",
  2359 => x"86c887e3",
  2360 => x"ef49e0c0",
  2361 => x"a4c487ec",
  2362 => x"f0496a4a",
  2363 => x"caf187f3",
  2364 => x"c184cc87",
  2365 => x"abb7c883",
  2366 => x"87cdff04",
  2367 => x"4d268efc",
  2368 => x"4b264c26",
  2369 => x"711e4f26",
  2370 => x"d8fcc24a",
  2371 => x"d8fcc25a",
  2372 => x"4978c748",
  2373 => x"2687e1fe",
  2374 => x"1e731e4f",
  2375 => x"b7c04a71",
  2376 => x"87d303aa",
  2377 => x"bffce0c2",
  2378 => x"c187c405",
  2379 => x"c087c24b",
  2380 => x"c0e1c24b",
  2381 => x"c287c45b",
  2382 => x"fc5ac0e1",
  2383 => x"fce0c248",
  2384 => x"c14a78bf",
  2385 => x"a2c0c19a",
  2386 => x"87e8ec49",
  2387 => x"4f264b26",
  2388 => x"c44a711e",
  2389 => x"49721e66",
  2390 => x"fc87e0eb",
  2391 => x"1e4f268e",
  2392 => x"c348d4ff",
  2393 => x"d0ff78ff",
  2394 => x"78e1c048",
  2395 => x"c148d4ff",
  2396 => x"c4487178",
  2397 => x"08d4ff30",
  2398 => x"48d0ff78",
  2399 => x"2678e0c0",
  2400 => x"5b5e0e4f",
  2401 => x"f00e5d5c",
  2402 => x"48a6c886",
  2403 => x"ec4d78c0",
  2404 => x"80fc7ebf",
  2405 => x"bfd4fcc2",
  2406 => x"4cbfe878",
  2407 => x"bffce0c2",
  2408 => x"87dde349",
  2409 => x"ca49eecb",
  2410 => x"4b7087d6",
  2411 => x"d2e749c7",
  2412 => x"05987087",
  2413 => x"496e87c8",
  2414 => x"c10299c1",
  2415 => x"4dc187c1",
  2416 => x"c27ebfec",
  2417 => x"49bffce0",
  2418 => x"7387f6e2",
  2419 => x"87fcc949",
  2420 => x"d7029870",
  2421 => x"f4e0c287",
  2422 => x"b9c149bf",
  2423 => x"59f8e0c2",
  2424 => x"87fbfd71",
  2425 => x"c949eecb",
  2426 => x"4b7087d6",
  2427 => x"d2e649c7",
  2428 => x"05987087",
  2429 => x"6e87c7ff",
  2430 => x"0599c149",
  2431 => x"7587fffe",
  2432 => x"e3c0029d",
  2433 => x"fce0c287",
  2434 => x"bac14abf",
  2435 => x"5ac0e1c2",
  2436 => x"0a7a0afc",
  2437 => x"c0c19ac1",
  2438 => x"d7e949a2",
  2439 => x"49dac187",
  2440 => x"c887e0e5",
  2441 => x"78c148a6",
  2442 => x"bffce0c2",
  2443 => x"87e9c005",
  2444 => x"ffc34974",
  2445 => x"c01e7199",
  2446 => x"87d4fc49",
  2447 => x"b7c84974",
  2448 => x"c11e7129",
  2449 => x"87c8fc49",
  2450 => x"fdc386c8",
  2451 => x"87f3e449",
  2452 => x"e449fac3",
  2453 => x"d1c787ed",
  2454 => x"c3497487",
  2455 => x"b7c899ff",
  2456 => x"74b4712c",
  2457 => x"87df029c",
  2458 => x"bff8e0c2",
  2459 => x"87dcc749",
  2460 => x"c0059870",
  2461 => x"4cc087c4",
  2462 => x"e0c287d3",
  2463 => x"87c0c749",
  2464 => x"58fce0c2",
  2465 => x"c287c6c0",
  2466 => x"c048f8e0",
  2467 => x"c8497478",
  2468 => x"87ce0599",
  2469 => x"e349f5c3",
  2470 => x"497087e9",
  2471 => x"c00299c2",
  2472 => x"fcc287e9",
  2473 => x"c002bfd8",
  2474 => x"c14887c9",
  2475 => x"dcfcc288",
  2476 => x"c487d358",
  2477 => x"e0c14866",
  2478 => x"6e7e7080",
  2479 => x"c5c002bf",
  2480 => x"49ff4b87",
  2481 => x"a6c80f73",
  2482 => x"7478c148",
  2483 => x"0599c449",
  2484 => x"c387cec0",
  2485 => x"eae249f2",
  2486 => x"c2497087",
  2487 => x"f0c00299",
  2488 => x"d8fcc287",
  2489 => x"c7487ebf",
  2490 => x"c003a8b7",
  2491 => x"486e87cb",
  2492 => x"fcc280c1",
  2493 => x"d3c058dc",
  2494 => x"4866c487",
  2495 => x"7080e0c1",
  2496 => x"02bf6e7e",
  2497 => x"4b87c5c0",
  2498 => x"0f7349fe",
  2499 => x"c148a6c8",
  2500 => x"49fdc378",
  2501 => x"7087ece1",
  2502 => x"0299c249",
  2503 => x"c287e9c0",
  2504 => x"02bfd8fc",
  2505 => x"c287c9c0",
  2506 => x"c048d8fc",
  2507 => x"87d3c078",
  2508 => x"c14866c4",
  2509 => x"7e7080e0",
  2510 => x"c002bf6e",
  2511 => x"fd4b87c5",
  2512 => x"c80f7349",
  2513 => x"78c148a6",
  2514 => x"e049fac3",
  2515 => x"497087f5",
  2516 => x"c00299c2",
  2517 => x"fcc287ea",
  2518 => x"c748bfd8",
  2519 => x"c003a8b7",
  2520 => x"fcc287c9",
  2521 => x"78c748d8",
  2522 => x"c487d0c0",
  2523 => x"e0c14a66",
  2524 => x"c0026a82",
  2525 => x"fc4b87c5",
  2526 => x"c80f7349",
  2527 => x"78c148a6",
  2528 => x"fcc24dc0",
  2529 => x"50c048d0",
  2530 => x"c249eecb",
  2531 => x"4b7087f2",
  2532 => x"97d0fcc2",
  2533 => x"ddc105bf",
  2534 => x"c3497487",
  2535 => x"c00599f0",
  2536 => x"dac187cd",
  2537 => x"dadfff49",
  2538 => x"02987087",
  2539 => x"c187c7c1",
  2540 => x"4cbfe84d",
  2541 => x"99ffc349",
  2542 => x"712cb7c8",
  2543 => x"fce0c2b4",
  2544 => x"daff49bf",
  2545 => x"497387fb",
  2546 => x"7087c1c2",
  2547 => x"c6c00298",
  2548 => x"d0fcc287",
  2549 => x"c250c148",
  2550 => x"bf97d0fc",
  2551 => x"87d6c005",
  2552 => x"f0c34974",
  2553 => x"c6ff0599",
  2554 => x"49dac187",
  2555 => x"87d3deff",
  2556 => x"fe059870",
  2557 => x"9d7587f9",
  2558 => x"87e0c002",
  2559 => x"c248a6cc",
  2560 => x"78bfd8fc",
  2561 => x"cc4966cc",
  2562 => x"4866c491",
  2563 => x"7e708071",
  2564 => x"c002bf6e",
  2565 => x"cc4b87c6",
  2566 => x"0f734966",
  2567 => x"c00266c8",
  2568 => x"fcc287c8",
  2569 => x"f249bfd8",
  2570 => x"8ef087ce",
  2571 => x"4c264d26",
  2572 => x"4f264b26",
  2573 => x"00000000",
  2574 => x"00000000",
  2575 => x"00000000",
  2576 => x"ff4a711e",
  2577 => x"7249bfc8",
  2578 => x"4f2648a1",
  2579 => x"bfc8ff1e",
  2580 => x"c0c0fe89",
  2581 => x"a9c0c0c0",
  2582 => x"c087c401",
  2583 => x"c187c24a",
  2584 => x"2648724a",
  2585 => x"5b5e0e4f",
  2586 => x"710e5d5c",
  2587 => x"4cd4ff4b",
  2588 => x"c04866d0",
  2589 => x"ff49d678",
  2590 => x"c387c5de",
  2591 => x"496c7cff",
  2592 => x"7199ffc3",
  2593 => x"f0c3494d",
  2594 => x"a9e0c199",
  2595 => x"c387cb05",
  2596 => x"486c7cff",
  2597 => x"66d098c3",
  2598 => x"ffc37808",
  2599 => x"494a6c7c",
  2600 => x"ffc331c8",
  2601 => x"714a6c7c",
  2602 => x"c84972b2",
  2603 => x"7cffc331",
  2604 => x"b2714a6c",
  2605 => x"31c84972",
  2606 => x"6c7cffc3",
  2607 => x"ffb2714a",
  2608 => x"e0c048d0",
  2609 => x"029b7378",
  2610 => x"7b7287c2",
  2611 => x"4d264875",
  2612 => x"4b264c26",
  2613 => x"261e4f26",
  2614 => x"5b5e0e4f",
  2615 => x"86f80e5c",
  2616 => x"a6c81e76",
  2617 => x"87fdfd49",
  2618 => x"4b7086c4",
  2619 => x"a8c4486e",
  2620 => x"87f4c203",
  2621 => x"f0c34a73",
  2622 => x"aad0c19a",
  2623 => x"c187c702",
  2624 => x"c205aae0",
  2625 => x"497387e2",
  2626 => x"c30299c8",
  2627 => x"87c6ff87",
  2628 => x"9cc34c73",
  2629 => x"c105acc2",
  2630 => x"66c487c4",
  2631 => x"7131c949",
  2632 => x"4a66c41e",
  2633 => x"c292c8c1",
  2634 => x"7249dcfc",
  2635 => x"c0ccfe81",
  2636 => x"ff49d887",
  2637 => x"c887c9db",
  2638 => x"eac21ec0",
  2639 => x"e1fd49c0",
  2640 => x"d0ff87fa",
  2641 => x"78e0c048",
  2642 => x"1ec0eac2",
  2643 => x"c14a66cc",
  2644 => x"fcc292c8",
  2645 => x"817249dc",
  2646 => x"87cac7fe",
  2647 => x"acc186cc",
  2648 => x"87c4c105",
  2649 => x"c94966c4",
  2650 => x"c41e7131",
  2651 => x"c8c14a66",
  2652 => x"dcfcc292",
  2653 => x"fe817249",
  2654 => x"c287f6ca",
  2655 => x"c81ec0ea",
  2656 => x"c8c14a66",
  2657 => x"dcfcc292",
  2658 => x"fe817249",
  2659 => x"d787c8c5",
  2660 => x"ebd9ff49",
  2661 => x"1ec0c887",
  2662 => x"49c0eac2",
  2663 => x"87f9dffd",
  2664 => x"d0ff86cc",
  2665 => x"78e0c048",
  2666 => x"4c268ef8",
  2667 => x"4f264b26",
  2668 => x"5c5b5e0e",
  2669 => x"86fc0e5d",
  2670 => x"d4ff4d71",
  2671 => x"7e66d44c",
  2672 => x"a8b7c348",
  2673 => x"87e3c101",
  2674 => x"66c41e75",
  2675 => x"93c8c14b",
  2676 => x"83dcfcc2",
  2677 => x"fdfd4973",
  2678 => x"a3c887ff",
  2679 => x"ff496949",
  2680 => x"e1c848d0",
  2681 => x"717cdd78",
  2682 => x"98ffc348",
  2683 => x"4a717c70",
  2684 => x"722ab7c8",
  2685 => x"98ffc348",
  2686 => x"4a717c70",
  2687 => x"722ab7d0",
  2688 => x"98ffc348",
  2689 => x"48717c70",
  2690 => x"7028b7d8",
  2691 => x"7c7cc07c",
  2692 => x"7c7c7c7c",
  2693 => x"7c7c7c7c",
  2694 => x"d0ff7c7c",
  2695 => x"78e0c048",
  2696 => x"dc1e66c4",
  2697 => x"fcd7ff49",
  2698 => x"fc86c887",
  2699 => x"264d268e",
  2700 => x"264b264c",
  2701 => x"e9c21e4f",
  2702 => x"fe49bfc4",
  2703 => x"c087efdc",
  2704 => x"004f2648",
  2705 => x"00002a48",
  2706 => x"54534d41",
  2707 => x"20444152",
  2708 => x"004d4f52",
  2709 => x"00001d97",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
